VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO leorv32
  CLASS BLOCK ;
  FOREIGN leorv32 ;
  ORIGIN 0.000 0.000 ;
  SIZE 500.000 BY 500.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.490 0.000 41.770 4.000 ;
    END
  END clk
  PIN mem_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.350 496.000 14.630 500.000 ;
    END
  END mem_addr[0]
  PIN mem_addr[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 166.150 496.000 166.430 500.000 ;
    END
  END mem_addr[10]
  PIN mem_addr[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 181.330 496.000 181.610 500.000 ;
    END
  END mem_addr[11]
  PIN mem_addr[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.510 496.000 196.790 500.000 ;
    END
  END mem_addr[12]
  PIN mem_addr[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 211.690 496.000 211.970 500.000 ;
    END
  END mem_addr[13]
  PIN mem_addr[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 226.870 496.000 227.150 500.000 ;
    END
  END mem_addr[14]
  PIN mem_addr[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.050 496.000 242.330 500.000 ;
    END
  END mem_addr[15]
  PIN mem_addr[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.230 496.000 257.510 500.000 ;
    END
  END mem_addr[16]
  PIN mem_addr[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 272.410 496.000 272.690 500.000 ;
    END
  END mem_addr[17]
  PIN mem_addr[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 287.590 496.000 287.870 500.000 ;
    END
  END mem_addr[18]
  PIN mem_addr[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.770 496.000 303.050 500.000 ;
    END
  END mem_addr[19]
  PIN mem_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.530 496.000 29.810 500.000 ;
    END
  END mem_addr[1]
  PIN mem_addr[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.950 496.000 318.230 500.000 ;
    END
  END mem_addr[20]
  PIN mem_addr[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 333.130 496.000 333.410 500.000 ;
    END
  END mem_addr[21]
  PIN mem_addr[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 348.310 496.000 348.590 500.000 ;
    END
  END mem_addr[22]
  PIN mem_addr[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.490 496.000 363.770 500.000 ;
    END
  END mem_addr[23]
  PIN mem_addr[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 378.670 496.000 378.950 500.000 ;
    END
  END mem_addr[24]
  PIN mem_addr[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 393.850 496.000 394.130 500.000 ;
    END
  END mem_addr[25]
  PIN mem_addr[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 409.030 496.000 409.310 500.000 ;
    END
  END mem_addr[26]
  PIN mem_addr[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 424.210 496.000 424.490 500.000 ;
    END
  END mem_addr[27]
  PIN mem_addr[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 439.390 496.000 439.670 500.000 ;
    END
  END mem_addr[28]
  PIN mem_addr[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 454.570 496.000 454.850 500.000 ;
    END
  END mem_addr[29]
  PIN mem_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.710 496.000 44.990 500.000 ;
    END
  END mem_addr[2]
  PIN mem_addr[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 469.750 496.000 470.030 500.000 ;
    END
  END mem_addr[30]
  PIN mem_addr[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 484.930 496.000 485.210 500.000 ;
    END
  END mem_addr[31]
  PIN mem_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.890 496.000 60.170 500.000 ;
    END
  END mem_addr[3]
  PIN mem_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.070 496.000 75.350 500.000 ;
    END
  END mem_addr[4]
  PIN mem_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.250 496.000 90.530 500.000 ;
    END
  END mem_addr[5]
  PIN mem_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.430 496.000 105.710 500.000 ;
    END
  END mem_addr[6]
  PIN mem_addr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.610 496.000 120.890 500.000 ;
    END
  END mem_addr[7]
  PIN mem_addr[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.790 496.000 136.070 500.000 ;
    END
  END mem_addr[8]
  PIN mem_addr[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.970 496.000 151.250 500.000 ;
    END
  END mem_addr[9]
  PIN mem_rbusy
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.530 0.000 374.810 4.000 ;
    END
  END mem_rbusy
  PIN mem_rdata[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.720 4.000 18.320 ;
    END
  END mem_rdata[0]
  PIN mem_rdata[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 167.320 4.000 167.920 ;
    END
  END mem_rdata[10]
  PIN mem_rdata[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 182.280 4.000 182.880 ;
    END
  END mem_rdata[11]
  PIN mem_rdata[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 197.240 4.000 197.840 ;
    END
  END mem_rdata[12]
  PIN mem_rdata[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 212.200 4.000 212.800 ;
    END
  END mem_rdata[13]
  PIN mem_rdata[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 227.160 4.000 227.760 ;
    END
  END mem_rdata[14]
  PIN mem_rdata[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 242.120 4.000 242.720 ;
    END
  END mem_rdata[15]
  PIN mem_rdata[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 257.080 4.000 257.680 ;
    END
  END mem_rdata[16]
  PIN mem_rdata[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 272.040 4.000 272.640 ;
    END
  END mem_rdata[17]
  PIN mem_rdata[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 287.000 4.000 287.600 ;
    END
  END mem_rdata[18]
  PIN mem_rdata[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 301.960 4.000 302.560 ;
    END
  END mem_rdata[19]
  PIN mem_rdata[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 32.680 4.000 33.280 ;
    END
  END mem_rdata[1]
  PIN mem_rdata[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 316.920 4.000 317.520 ;
    END
  END mem_rdata[20]
  PIN mem_rdata[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 331.880 4.000 332.480 ;
    END
  END mem_rdata[21]
  PIN mem_rdata[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 346.840 4.000 347.440 ;
    END
  END mem_rdata[22]
  PIN mem_rdata[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 361.800 4.000 362.400 ;
    END
  END mem_rdata[23]
  PIN mem_rdata[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 376.760 4.000 377.360 ;
    END
  END mem_rdata[24]
  PIN mem_rdata[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 391.720 4.000 392.320 ;
    END
  END mem_rdata[25]
  PIN mem_rdata[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 406.680 4.000 407.280 ;
    END
  END mem_rdata[26]
  PIN mem_rdata[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 421.640 4.000 422.240 ;
    END
  END mem_rdata[27]
  PIN mem_rdata[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 436.600 4.000 437.200 ;
    END
  END mem_rdata[28]
  PIN mem_rdata[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 451.560 4.000 452.160 ;
    END
  END mem_rdata[29]
  PIN mem_rdata[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 4.000 48.240 ;
    END
  END mem_rdata[2]
  PIN mem_rdata[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 466.520 4.000 467.120 ;
    END
  END mem_rdata[30]
  PIN mem_rdata[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 481.480 4.000 482.080 ;
    END
  END mem_rdata[31]
  PIN mem_rdata[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 62.600 4.000 63.200 ;
    END
  END mem_rdata[3]
  PIN mem_rdata[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 77.560 4.000 78.160 ;
    END
  END mem_rdata[4]
  PIN mem_rdata[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 92.520 4.000 93.120 ;
    END
  END mem_rdata[5]
  PIN mem_rdata[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 107.480 4.000 108.080 ;
    END
  END mem_rdata[6]
  PIN mem_rdata[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 122.440 4.000 123.040 ;
    END
  END mem_rdata[7]
  PIN mem_rdata[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 137.400 4.000 138.000 ;
    END
  END mem_rdata[8]
  PIN mem_rdata[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 152.360 4.000 152.960 ;
    END
  END mem_rdata[9]
  PIN mem_rstrb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 291.270 0.000 291.550 4.000 ;
    END
  END mem_rstrb
  PIN mem_wbusy
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 457.790 0.000 458.070 4.000 ;
    END
  END mem_wbusy
  PIN mem_wdata[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 11.600 500.000 12.200 ;
    END
  END mem_wdata[0]
  PIN mem_wdata[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 147.600 500.000 148.200 ;
    END
  END mem_wdata[10]
  PIN mem_wdata[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 161.200 500.000 161.800 ;
    END
  END mem_wdata[11]
  PIN mem_wdata[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 174.800 500.000 175.400 ;
    END
  END mem_wdata[12]
  PIN mem_wdata[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 188.400 500.000 189.000 ;
    END
  END mem_wdata[13]
  PIN mem_wdata[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 202.000 500.000 202.600 ;
    END
  END mem_wdata[14]
  PIN mem_wdata[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 215.600 500.000 216.200 ;
    END
  END mem_wdata[15]
  PIN mem_wdata[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 229.200 500.000 229.800 ;
    END
  END mem_wdata[16]
  PIN mem_wdata[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 242.800 500.000 243.400 ;
    END
  END mem_wdata[17]
  PIN mem_wdata[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 256.400 500.000 257.000 ;
    END
  END mem_wdata[18]
  PIN mem_wdata[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 270.000 500.000 270.600 ;
    END
  END mem_wdata[19]
  PIN mem_wdata[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 25.200 500.000 25.800 ;
    END
  END mem_wdata[1]
  PIN mem_wdata[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 283.600 500.000 284.200 ;
    END
  END mem_wdata[20]
  PIN mem_wdata[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 297.200 500.000 297.800 ;
    END
  END mem_wdata[21]
  PIN mem_wdata[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 310.800 500.000 311.400 ;
    END
  END mem_wdata[22]
  PIN mem_wdata[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 324.400 500.000 325.000 ;
    END
  END mem_wdata[23]
  PIN mem_wdata[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 338.000 500.000 338.600 ;
    END
  END mem_wdata[24]
  PIN mem_wdata[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 351.600 500.000 352.200 ;
    END
  END mem_wdata[25]
  PIN mem_wdata[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 365.200 500.000 365.800 ;
    END
  END mem_wdata[26]
  PIN mem_wdata[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 378.800 500.000 379.400 ;
    END
  END mem_wdata[27]
  PIN mem_wdata[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 392.400 500.000 393.000 ;
    END
  END mem_wdata[28]
  PIN mem_wdata[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 406.000 500.000 406.600 ;
    END
  END mem_wdata[29]
  PIN mem_wdata[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 38.800 500.000 39.400 ;
    END
  END mem_wdata[2]
  PIN mem_wdata[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 419.600 500.000 420.200 ;
    END
  END mem_wdata[30]
  PIN mem_wdata[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 433.200 500.000 433.800 ;
    END
  END mem_wdata[31]
  PIN mem_wdata[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 52.400 500.000 53.000 ;
    END
  END mem_wdata[3]
  PIN mem_wdata[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 66.000 500.000 66.600 ;
    END
  END mem_wdata[4]
  PIN mem_wdata[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 79.600 500.000 80.200 ;
    END
  END mem_wdata[5]
  PIN mem_wdata[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 93.200 500.000 93.800 ;
    END
  END mem_wdata[6]
  PIN mem_wdata[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 106.800 500.000 107.400 ;
    END
  END mem_wdata[7]
  PIN mem_wdata[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 120.400 500.000 121.000 ;
    END
  END mem_wdata[8]
  PIN mem_wdata[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 134.000 500.000 134.600 ;
    END
  END mem_wdata[9]
  PIN mem_wmask[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 446.800 500.000 447.400 ;
    END
  END mem_wmask[0]
  PIN mem_wmask[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 460.400 500.000 461.000 ;
    END
  END mem_wmask[1]
  PIN mem_wmask[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 474.000 500.000 474.600 ;
    END
  END mem_wmask[2]
  PIN mem_wmask[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 487.600 500.000 488.200 ;
    END
  END mem_wmask[3]
  PIN mhartid_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.010 0.000 208.290 4.000 ;
    END
  END mhartid_0
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.750 0.000 125.030 4.000 ;
    END
  END reset
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 487.120 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 487.120 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 494.040 486.965 ;
      LAYER met1 ;
        RECT 1.450 2.080 499.950 489.560 ;
      LAYER met2 ;
        RECT 0.090 495.720 14.070 496.810 ;
        RECT 14.910 495.720 29.250 496.810 ;
        RECT 30.090 495.720 44.430 496.810 ;
        RECT 45.270 495.720 59.610 496.810 ;
        RECT 60.450 495.720 74.790 496.810 ;
        RECT 75.630 495.720 89.970 496.810 ;
        RECT 90.810 495.720 105.150 496.810 ;
        RECT 105.990 495.720 120.330 496.810 ;
        RECT 121.170 495.720 135.510 496.810 ;
        RECT 136.350 495.720 150.690 496.810 ;
        RECT 151.530 495.720 165.870 496.810 ;
        RECT 166.710 495.720 181.050 496.810 ;
        RECT 181.890 495.720 196.230 496.810 ;
        RECT 197.070 495.720 211.410 496.810 ;
        RECT 212.250 495.720 226.590 496.810 ;
        RECT 227.430 495.720 241.770 496.810 ;
        RECT 242.610 495.720 256.950 496.810 ;
        RECT 257.790 495.720 272.130 496.810 ;
        RECT 272.970 495.720 287.310 496.810 ;
        RECT 288.150 495.720 302.490 496.810 ;
        RECT 303.330 495.720 317.670 496.810 ;
        RECT 318.510 495.720 332.850 496.810 ;
        RECT 333.690 495.720 348.030 496.810 ;
        RECT 348.870 495.720 363.210 496.810 ;
        RECT 364.050 495.720 378.390 496.810 ;
        RECT 379.230 495.720 393.570 496.810 ;
        RECT 394.410 495.720 408.750 496.810 ;
        RECT 409.590 495.720 423.930 496.810 ;
        RECT 424.770 495.720 439.110 496.810 ;
        RECT 439.950 495.720 454.290 496.810 ;
        RECT 455.130 495.720 469.470 496.810 ;
        RECT 470.310 495.720 484.650 496.810 ;
        RECT 485.490 495.720 499.920 496.810 ;
        RECT 0.090 4.280 499.920 495.720 ;
        RECT 0.090 0.155 41.210 4.280 ;
        RECT 42.050 0.155 124.470 4.280 ;
        RECT 125.310 0.155 207.730 4.280 ;
        RECT 208.570 0.155 290.990 4.280 ;
        RECT 291.830 0.155 374.250 4.280 ;
        RECT 375.090 0.155 457.510 4.280 ;
        RECT 458.350 0.155 499.920 4.280 ;
      LAYER met3 ;
        RECT 0.065 487.200 495.600 488.065 ;
        RECT 0.065 482.480 499.495 487.200 ;
        RECT 4.400 481.080 499.495 482.480 ;
        RECT 0.065 475.000 499.495 481.080 ;
        RECT 0.065 473.600 495.600 475.000 ;
        RECT 0.065 467.520 499.495 473.600 ;
        RECT 4.400 466.120 499.495 467.520 ;
        RECT 0.065 461.400 499.495 466.120 ;
        RECT 0.065 460.000 495.600 461.400 ;
        RECT 0.065 452.560 499.495 460.000 ;
        RECT 4.400 451.160 499.495 452.560 ;
        RECT 0.065 447.800 499.495 451.160 ;
        RECT 0.065 446.400 495.600 447.800 ;
        RECT 0.065 437.600 499.495 446.400 ;
        RECT 4.400 436.200 499.495 437.600 ;
        RECT 0.065 434.200 499.495 436.200 ;
        RECT 0.065 432.800 495.600 434.200 ;
        RECT 0.065 422.640 499.495 432.800 ;
        RECT 4.400 421.240 499.495 422.640 ;
        RECT 0.065 420.600 499.495 421.240 ;
        RECT 0.065 419.200 495.600 420.600 ;
        RECT 0.065 407.680 499.495 419.200 ;
        RECT 4.400 407.000 499.495 407.680 ;
        RECT 4.400 406.280 495.600 407.000 ;
        RECT 0.065 405.600 495.600 406.280 ;
        RECT 0.065 393.400 499.495 405.600 ;
        RECT 0.065 392.720 495.600 393.400 ;
        RECT 4.400 392.000 495.600 392.720 ;
        RECT 4.400 391.320 499.495 392.000 ;
        RECT 0.065 379.800 499.495 391.320 ;
        RECT 0.065 378.400 495.600 379.800 ;
        RECT 0.065 377.760 499.495 378.400 ;
        RECT 4.400 376.360 499.495 377.760 ;
        RECT 0.065 366.200 499.495 376.360 ;
        RECT 0.065 364.800 495.600 366.200 ;
        RECT 0.065 362.800 499.495 364.800 ;
        RECT 4.400 361.400 499.495 362.800 ;
        RECT 0.065 352.600 499.495 361.400 ;
        RECT 0.065 351.200 495.600 352.600 ;
        RECT 0.065 347.840 499.495 351.200 ;
        RECT 4.400 346.440 499.495 347.840 ;
        RECT 0.065 339.000 499.495 346.440 ;
        RECT 0.065 337.600 495.600 339.000 ;
        RECT 0.065 332.880 499.495 337.600 ;
        RECT 4.400 331.480 499.495 332.880 ;
        RECT 0.065 325.400 499.495 331.480 ;
        RECT 0.065 324.000 495.600 325.400 ;
        RECT 0.065 317.920 499.495 324.000 ;
        RECT 4.400 316.520 499.495 317.920 ;
        RECT 0.065 311.800 499.495 316.520 ;
        RECT 0.065 310.400 495.600 311.800 ;
        RECT 0.065 302.960 499.495 310.400 ;
        RECT 4.400 301.560 499.495 302.960 ;
        RECT 0.065 298.200 499.495 301.560 ;
        RECT 0.065 296.800 495.600 298.200 ;
        RECT 0.065 288.000 499.495 296.800 ;
        RECT 4.400 286.600 499.495 288.000 ;
        RECT 0.065 284.600 499.495 286.600 ;
        RECT 0.065 283.200 495.600 284.600 ;
        RECT 0.065 273.040 499.495 283.200 ;
        RECT 4.400 271.640 499.495 273.040 ;
        RECT 0.065 271.000 499.495 271.640 ;
        RECT 0.065 269.600 495.600 271.000 ;
        RECT 0.065 258.080 499.495 269.600 ;
        RECT 4.400 257.400 499.495 258.080 ;
        RECT 4.400 256.680 495.600 257.400 ;
        RECT 0.065 256.000 495.600 256.680 ;
        RECT 0.065 243.800 499.495 256.000 ;
        RECT 0.065 243.120 495.600 243.800 ;
        RECT 4.400 242.400 495.600 243.120 ;
        RECT 4.400 241.720 499.495 242.400 ;
        RECT 0.065 230.200 499.495 241.720 ;
        RECT 0.065 228.800 495.600 230.200 ;
        RECT 0.065 228.160 499.495 228.800 ;
        RECT 4.400 226.760 499.495 228.160 ;
        RECT 0.065 216.600 499.495 226.760 ;
        RECT 0.065 215.200 495.600 216.600 ;
        RECT 0.065 213.200 499.495 215.200 ;
        RECT 4.400 211.800 499.495 213.200 ;
        RECT 0.065 203.000 499.495 211.800 ;
        RECT 0.065 201.600 495.600 203.000 ;
        RECT 0.065 198.240 499.495 201.600 ;
        RECT 4.400 196.840 499.495 198.240 ;
        RECT 0.065 189.400 499.495 196.840 ;
        RECT 0.065 188.000 495.600 189.400 ;
        RECT 0.065 183.280 499.495 188.000 ;
        RECT 4.400 181.880 499.495 183.280 ;
        RECT 0.065 175.800 499.495 181.880 ;
        RECT 0.065 174.400 495.600 175.800 ;
        RECT 0.065 168.320 499.495 174.400 ;
        RECT 4.400 166.920 499.495 168.320 ;
        RECT 0.065 162.200 499.495 166.920 ;
        RECT 0.065 160.800 495.600 162.200 ;
        RECT 0.065 153.360 499.495 160.800 ;
        RECT 4.400 151.960 499.495 153.360 ;
        RECT 0.065 148.600 499.495 151.960 ;
        RECT 0.065 147.200 495.600 148.600 ;
        RECT 0.065 138.400 499.495 147.200 ;
        RECT 4.400 137.000 499.495 138.400 ;
        RECT 0.065 135.000 499.495 137.000 ;
        RECT 0.065 133.600 495.600 135.000 ;
        RECT 0.065 123.440 499.495 133.600 ;
        RECT 4.400 122.040 499.495 123.440 ;
        RECT 0.065 121.400 499.495 122.040 ;
        RECT 0.065 120.000 495.600 121.400 ;
        RECT 0.065 108.480 499.495 120.000 ;
        RECT 4.400 107.800 499.495 108.480 ;
        RECT 4.400 107.080 495.600 107.800 ;
        RECT 0.065 106.400 495.600 107.080 ;
        RECT 0.065 94.200 499.495 106.400 ;
        RECT 0.065 93.520 495.600 94.200 ;
        RECT 4.400 92.800 495.600 93.520 ;
        RECT 4.400 92.120 499.495 92.800 ;
        RECT 0.065 80.600 499.495 92.120 ;
        RECT 0.065 79.200 495.600 80.600 ;
        RECT 0.065 78.560 499.495 79.200 ;
        RECT 4.400 77.160 499.495 78.560 ;
        RECT 0.065 67.000 499.495 77.160 ;
        RECT 0.065 65.600 495.600 67.000 ;
        RECT 0.065 63.600 499.495 65.600 ;
        RECT 4.400 62.200 499.495 63.600 ;
        RECT 0.065 53.400 499.495 62.200 ;
        RECT 0.065 52.000 495.600 53.400 ;
        RECT 0.065 48.640 499.495 52.000 ;
        RECT 4.400 47.240 499.495 48.640 ;
        RECT 0.065 39.800 499.495 47.240 ;
        RECT 0.065 38.400 495.600 39.800 ;
        RECT 0.065 33.680 499.495 38.400 ;
        RECT 4.400 32.280 499.495 33.680 ;
        RECT 0.065 26.200 499.495 32.280 ;
        RECT 0.065 24.800 495.600 26.200 ;
        RECT 0.065 18.720 499.495 24.800 ;
        RECT 4.400 17.320 499.495 18.720 ;
        RECT 0.065 12.600 499.495 17.320 ;
        RECT 0.065 11.200 495.600 12.600 ;
        RECT 0.065 0.175 499.495 11.200 ;
      LAYER met4 ;
        RECT 2.135 10.240 20.640 486.025 ;
        RECT 23.040 10.240 97.440 486.025 ;
        RECT 99.840 10.240 174.240 486.025 ;
        RECT 176.640 10.240 251.040 486.025 ;
        RECT 253.440 10.240 327.840 486.025 ;
        RECT 330.240 10.240 404.640 486.025 ;
        RECT 407.040 10.240 481.440 486.025 ;
        RECT 483.840 10.240 499.265 486.025 ;
        RECT 2.135 0.175 499.265 10.240 ;
  END
END leorv32
END LIBRARY

