// This is the unpowered netlist.
module leorv32 (clk,
    mem_rbusy,
    mem_rstrb,
    mem_wbusy,
    mhartid_0,
    reset,
    mem_addr,
    mem_rdata,
    mem_wdata,
    mem_wmask);
 input clk;
 input mem_rbusy;
 output mem_rstrb;
 input mem_wbusy;
 input mhartid_0;
 input reset;
 output [31:0] mem_addr;
 input [31:0] mem_rdata;
 output [31:0] mem_wdata;
 output [3:0] mem_wmask;

 wire \B_type_imm[11] ;
 wire \B_type_imm[12] ;
 wire \B_type_imm[1] ;
 wire \B_type_imm[2] ;
 wire \B_type_imm[3] ;
 wire \B_type_imm[4] ;
 wire \B_type_imm[5] ;
 wire \B_type_imm[6] ;
 wire \B_type_imm[7] ;
 wire \B_type_imm[8] ;
 wire \B_type_imm[9] ;
 wire \I_type_imm[0] ;
 wire \I_type_imm[1] ;
 wire \I_type_imm[2] ;
 wire \I_type_imm[3] ;
 wire \I_type_imm[4] ;
 wire \J_type_imm[12] ;
 wire \J_type_imm[13] ;
 wire \J_type_imm[14] ;
 wire \J_type_imm[15] ;
 wire \J_type_imm[16] ;
 wire \J_type_imm[17] ;
 wire \J_type_imm[18] ;
 wire \J_type_imm[19] ;
 wire \PC[10] ;
 wire \PC[11] ;
 wire \PC[12] ;
 wire \PC[13] ;
 wire \PC[14] ;
 wire \PC[15] ;
 wire \PC[16] ;
 wire \PC[17] ;
 wire \PC[18] ;
 wire \PC[19] ;
 wire \PC[1] ;
 wire \PC[20] ;
 wire \PC[21] ;
 wire \PC[22] ;
 wire \PC[23] ;
 wire \PC[2] ;
 wire \PC[3] ;
 wire \PC[4] ;
 wire \PC[5] ;
 wire \PC[6] ;
 wire \PC[7] ;
 wire \PC[8] ;
 wire \PC[9] ;
 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire _06906_;
 wire _06907_;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire _06911_;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire _06921_;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire _06928_;
 wire _06929_;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire _06937_;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire _06948_;
 wire _06949_;
 wire _06950_;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire _06965_;
 wire _06966_;
 wire _06967_;
 wire _06968_;
 wire _06969_;
 wire _06970_;
 wire _06971_;
 wire _06972_;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire _06976_;
 wire _06977_;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire _06982_;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire _06987_;
 wire _06988_;
 wire _06989_;
 wire _06990_;
 wire _06991_;
 wire _06992_;
 wire _06993_;
 wire _06994_;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire _07000_;
 wire _07001_;
 wire _07002_;
 wire _07003_;
 wire _07004_;
 wire _07005_;
 wire _07006_;
 wire _07007_;
 wire _07008_;
 wire _07009_;
 wire _07010_;
 wire _07011_;
 wire _07012_;
 wire _07013_;
 wire _07014_;
 wire _07015_;
 wire _07016_;
 wire _07017_;
 wire _07018_;
 wire _07019_;
 wire _07020_;
 wire _07021_;
 wire _07022_;
 wire _07023_;
 wire _07024_;
 wire _07025_;
 wire _07026_;
 wire _07027_;
 wire _07028_;
 wire _07029_;
 wire _07030_;
 wire _07031_;
 wire \barrel_shifter_right.arith ;
 wire \core_state[0] ;
 wire \core_state[1] ;
 wire \core_state[2] ;
 wire \core_state[3] ;
 wire \cycles[0] ;
 wire \cycles[10] ;
 wire \cycles[11] ;
 wire \cycles[12] ;
 wire \cycles[13] ;
 wire \cycles[14] ;
 wire \cycles[15] ;
 wire \cycles[16] ;
 wire \cycles[17] ;
 wire \cycles[18] ;
 wire \cycles[19] ;
 wire \cycles[1] ;
 wire \cycles[20] ;
 wire \cycles[21] ;
 wire \cycles[22] ;
 wire \cycles[23] ;
 wire \cycles[24] ;
 wire \cycles[25] ;
 wire \cycles[26] ;
 wire \cycles[27] ;
 wire \cycles[28] ;
 wire \cycles[29] ;
 wire \cycles[2] ;
 wire \cycles[30] ;
 wire \cycles[31] ;
 wire \cycles[32] ;
 wire \cycles[33] ;
 wire \cycles[34] ;
 wire \cycles[35] ;
 wire \cycles[36] ;
 wire \cycles[37] ;
 wire \cycles[38] ;
 wire \cycles[39] ;
 wire \cycles[3] ;
 wire \cycles[40] ;
 wire \cycles[41] ;
 wire \cycles[42] ;
 wire \cycles[43] ;
 wire \cycles[44] ;
 wire \cycles[45] ;
 wire \cycles[46] ;
 wire \cycles[47] ;
 wire \cycles[48] ;
 wire \cycles[49] ;
 wire \cycles[4] ;
 wire \cycles[50] ;
 wire \cycles[51] ;
 wire \cycles[52] ;
 wire \cycles[53] ;
 wire \cycles[54] ;
 wire \cycles[55] ;
 wire \cycles[56] ;
 wire \cycles[57] ;
 wire \cycles[58] ;
 wire \cycles[59] ;
 wire \cycles[5] ;
 wire \cycles[60] ;
 wire \cycles[61] ;
 wire \cycles[62] ;
 wire \cycles[63] ;
 wire \cycles[6] ;
 wire \cycles[7] ;
 wire \cycles[8] ;
 wire \cycles[9] ;
 wire \instr[0] ;
 wire \instr[1] ;
 wire \instr[2] ;
 wire \instr[3] ;
 wire \instr[4] ;
 wire \instr[5] ;
 wire \instr[6] ;
 wire \instret[0] ;
 wire \instret[10] ;
 wire \instret[11] ;
 wire \instret[12] ;
 wire \instret[13] ;
 wire \instret[14] ;
 wire \instret[15] ;
 wire \instret[16] ;
 wire \instret[17] ;
 wire \instret[18] ;
 wire \instret[19] ;
 wire \instret[1] ;
 wire \instret[20] ;
 wire \instret[21] ;
 wire \instret[22] ;
 wire \instret[23] ;
 wire \instret[24] ;
 wire \instret[25] ;
 wire \instret[26] ;
 wire \instret[27] ;
 wire \instret[28] ;
 wire \instret[29] ;
 wire \instret[2] ;
 wire \instret[30] ;
 wire \instret[31] ;
 wire \instret[32] ;
 wire \instret[33] ;
 wire \instret[34] ;
 wire \instret[35] ;
 wire \instret[36] ;
 wire \instret[37] ;
 wire \instret[38] ;
 wire \instret[39] ;
 wire \instret[3] ;
 wire \instret[40] ;
 wire \instret[41] ;
 wire \instret[42] ;
 wire \instret[43] ;
 wire \instret[44] ;
 wire \instret[45] ;
 wire \instret[46] ;
 wire \instret[47] ;
 wire \instret[48] ;
 wire \instret[49] ;
 wire \instret[4] ;
 wire \instret[50] ;
 wire \instret[51] ;
 wire \instret[52] ;
 wire \instret[53] ;
 wire \instret[54] ;
 wire \instret[55] ;
 wire \instret[56] ;
 wire \instret[57] ;
 wire \instret[58] ;
 wire \instret[59] ;
 wire \instret[5] ;
 wire \instret[60] ;
 wire \instret[61] ;
 wire \instret[62] ;
 wire \instret[63] ;
 wire \instret[6] ;
 wire \instret[7] ;
 wire \instret[8] ;
 wire \instret[9] ;
 wire \leorv32_alu.input1[0] ;
 wire \leorv32_alu.input1[10] ;
 wire \leorv32_alu.input1[11] ;
 wire \leorv32_alu.input1[12] ;
 wire \leorv32_alu.input1[13] ;
 wire \leorv32_alu.input1[14] ;
 wire \leorv32_alu.input1[15] ;
 wire \leorv32_alu.input1[16] ;
 wire \leorv32_alu.input1[17] ;
 wire \leorv32_alu.input1[18] ;
 wire \leorv32_alu.input1[19] ;
 wire \leorv32_alu.input1[1] ;
 wire \leorv32_alu.input1[20] ;
 wire \leorv32_alu.input1[21] ;
 wire \leorv32_alu.input1[22] ;
 wire \leorv32_alu.input1[23] ;
 wire \leorv32_alu.input1[24] ;
 wire \leorv32_alu.input1[25] ;
 wire \leorv32_alu.input1[26] ;
 wire \leorv32_alu.input1[27] ;
 wire \leorv32_alu.input1[28] ;
 wire \leorv32_alu.input1[29] ;
 wire \leorv32_alu.input1[2] ;
 wire \leorv32_alu.input1[30] ;
 wire \leorv32_alu.input1[31] ;
 wire \leorv32_alu.input1[3] ;
 wire \leorv32_alu.input1[4] ;
 wire \leorv32_alu.input1[5] ;
 wire \leorv32_alu.input1[6] ;
 wire \leorv32_alu.input1[7] ;
 wire \leorv32_alu.input1[8] ;
 wire \leorv32_alu.input1[9] ;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire clknet_leaf_0_clk;
 wire \regs[0][0] ;
 wire \regs[0][10] ;
 wire \regs[0][11] ;
 wire \regs[0][12] ;
 wire \regs[0][13] ;
 wire \regs[0][14] ;
 wire \regs[0][15] ;
 wire \regs[0][16] ;
 wire \regs[0][17] ;
 wire \regs[0][18] ;
 wire \regs[0][19] ;
 wire \regs[0][1] ;
 wire \regs[0][20] ;
 wire \regs[0][21] ;
 wire \regs[0][22] ;
 wire \regs[0][23] ;
 wire \regs[0][24] ;
 wire \regs[0][25] ;
 wire \regs[0][26] ;
 wire \regs[0][27] ;
 wire \regs[0][28] ;
 wire \regs[0][29] ;
 wire \regs[0][2] ;
 wire \regs[0][30] ;
 wire \regs[0][31] ;
 wire \regs[0][3] ;
 wire \regs[0][4] ;
 wire \regs[0][5] ;
 wire \regs[0][6] ;
 wire \regs[0][7] ;
 wire \regs[0][8] ;
 wire \regs[0][9] ;
 wire \regs[10][0] ;
 wire \regs[10][10] ;
 wire \regs[10][11] ;
 wire \regs[10][12] ;
 wire \regs[10][13] ;
 wire \regs[10][14] ;
 wire \regs[10][15] ;
 wire \regs[10][16] ;
 wire \regs[10][17] ;
 wire \regs[10][18] ;
 wire \regs[10][19] ;
 wire \regs[10][1] ;
 wire \regs[10][20] ;
 wire \regs[10][21] ;
 wire \regs[10][22] ;
 wire \regs[10][23] ;
 wire \regs[10][24] ;
 wire \regs[10][25] ;
 wire \regs[10][26] ;
 wire \regs[10][27] ;
 wire \regs[10][28] ;
 wire \regs[10][29] ;
 wire \regs[10][2] ;
 wire \regs[10][30] ;
 wire \regs[10][31] ;
 wire \regs[10][3] ;
 wire \regs[10][4] ;
 wire \regs[10][5] ;
 wire \regs[10][6] ;
 wire \regs[10][7] ;
 wire \regs[10][8] ;
 wire \regs[10][9] ;
 wire \regs[11][0] ;
 wire \regs[11][10] ;
 wire \regs[11][11] ;
 wire \regs[11][12] ;
 wire \regs[11][13] ;
 wire \regs[11][14] ;
 wire \regs[11][15] ;
 wire \regs[11][16] ;
 wire \regs[11][17] ;
 wire \regs[11][18] ;
 wire \regs[11][19] ;
 wire \regs[11][1] ;
 wire \regs[11][20] ;
 wire \regs[11][21] ;
 wire \regs[11][22] ;
 wire \regs[11][23] ;
 wire \regs[11][24] ;
 wire \regs[11][25] ;
 wire \regs[11][26] ;
 wire \regs[11][27] ;
 wire \regs[11][28] ;
 wire \regs[11][29] ;
 wire \regs[11][2] ;
 wire \regs[11][30] ;
 wire \regs[11][31] ;
 wire \regs[11][3] ;
 wire \regs[11][4] ;
 wire \regs[11][5] ;
 wire \regs[11][6] ;
 wire \regs[11][7] ;
 wire \regs[11][8] ;
 wire \regs[11][9] ;
 wire \regs[12][0] ;
 wire \regs[12][10] ;
 wire \regs[12][11] ;
 wire \regs[12][12] ;
 wire \regs[12][13] ;
 wire \regs[12][14] ;
 wire \regs[12][15] ;
 wire \regs[12][16] ;
 wire \regs[12][17] ;
 wire \regs[12][18] ;
 wire \regs[12][19] ;
 wire \regs[12][1] ;
 wire \regs[12][20] ;
 wire \regs[12][21] ;
 wire \regs[12][22] ;
 wire \regs[12][23] ;
 wire \regs[12][24] ;
 wire \regs[12][25] ;
 wire \regs[12][26] ;
 wire \regs[12][27] ;
 wire \regs[12][28] ;
 wire \regs[12][29] ;
 wire \regs[12][2] ;
 wire \regs[12][30] ;
 wire \regs[12][31] ;
 wire \regs[12][3] ;
 wire \regs[12][4] ;
 wire \regs[12][5] ;
 wire \regs[12][6] ;
 wire \regs[12][7] ;
 wire \regs[12][8] ;
 wire \regs[12][9] ;
 wire \regs[13][0] ;
 wire \regs[13][10] ;
 wire \regs[13][11] ;
 wire \regs[13][12] ;
 wire \regs[13][13] ;
 wire \regs[13][14] ;
 wire \regs[13][15] ;
 wire \regs[13][16] ;
 wire \regs[13][17] ;
 wire \regs[13][18] ;
 wire \regs[13][19] ;
 wire \regs[13][1] ;
 wire \regs[13][20] ;
 wire \regs[13][21] ;
 wire \regs[13][22] ;
 wire \regs[13][23] ;
 wire \regs[13][24] ;
 wire \regs[13][25] ;
 wire \regs[13][26] ;
 wire \regs[13][27] ;
 wire \regs[13][28] ;
 wire \regs[13][29] ;
 wire \regs[13][2] ;
 wire \regs[13][30] ;
 wire \regs[13][31] ;
 wire \regs[13][3] ;
 wire \regs[13][4] ;
 wire \regs[13][5] ;
 wire \regs[13][6] ;
 wire \regs[13][7] ;
 wire \regs[13][8] ;
 wire \regs[13][9] ;
 wire \regs[14][0] ;
 wire \regs[14][10] ;
 wire \regs[14][11] ;
 wire \regs[14][12] ;
 wire \regs[14][13] ;
 wire \regs[14][14] ;
 wire \regs[14][15] ;
 wire \regs[14][16] ;
 wire \regs[14][17] ;
 wire \regs[14][18] ;
 wire \regs[14][19] ;
 wire \regs[14][1] ;
 wire \regs[14][20] ;
 wire \regs[14][21] ;
 wire \regs[14][22] ;
 wire \regs[14][23] ;
 wire \regs[14][24] ;
 wire \regs[14][25] ;
 wire \regs[14][26] ;
 wire \regs[14][27] ;
 wire \regs[14][28] ;
 wire \regs[14][29] ;
 wire \regs[14][2] ;
 wire \regs[14][30] ;
 wire \regs[14][31] ;
 wire \regs[14][3] ;
 wire \regs[14][4] ;
 wire \regs[14][5] ;
 wire \regs[14][6] ;
 wire \regs[14][7] ;
 wire \regs[14][8] ;
 wire \regs[14][9] ;
 wire \regs[15][0] ;
 wire \regs[15][10] ;
 wire \regs[15][11] ;
 wire \regs[15][12] ;
 wire \regs[15][13] ;
 wire \regs[15][14] ;
 wire \regs[15][15] ;
 wire \regs[15][16] ;
 wire \regs[15][17] ;
 wire \regs[15][18] ;
 wire \regs[15][19] ;
 wire \regs[15][1] ;
 wire \regs[15][20] ;
 wire \regs[15][21] ;
 wire \regs[15][22] ;
 wire \regs[15][23] ;
 wire \regs[15][24] ;
 wire \regs[15][25] ;
 wire \regs[15][26] ;
 wire \regs[15][27] ;
 wire \regs[15][28] ;
 wire \regs[15][29] ;
 wire \regs[15][2] ;
 wire \regs[15][30] ;
 wire \regs[15][31] ;
 wire \regs[15][3] ;
 wire \regs[15][4] ;
 wire \regs[15][5] ;
 wire \regs[15][6] ;
 wire \regs[15][7] ;
 wire \regs[15][8] ;
 wire \regs[15][9] ;
 wire \regs[16][0] ;
 wire \regs[16][10] ;
 wire \regs[16][11] ;
 wire \regs[16][12] ;
 wire \regs[16][13] ;
 wire \regs[16][14] ;
 wire \regs[16][15] ;
 wire \regs[16][16] ;
 wire \regs[16][17] ;
 wire \regs[16][18] ;
 wire \regs[16][19] ;
 wire \regs[16][1] ;
 wire \regs[16][20] ;
 wire \regs[16][21] ;
 wire \regs[16][22] ;
 wire \regs[16][23] ;
 wire \regs[16][24] ;
 wire \regs[16][25] ;
 wire \regs[16][26] ;
 wire \regs[16][27] ;
 wire \regs[16][28] ;
 wire \regs[16][29] ;
 wire \regs[16][2] ;
 wire \regs[16][30] ;
 wire \regs[16][31] ;
 wire \regs[16][3] ;
 wire \regs[16][4] ;
 wire \regs[16][5] ;
 wire \regs[16][6] ;
 wire \regs[16][7] ;
 wire \regs[16][8] ;
 wire \regs[16][9] ;
 wire \regs[17][0] ;
 wire \regs[17][10] ;
 wire \regs[17][11] ;
 wire \regs[17][12] ;
 wire \regs[17][13] ;
 wire \regs[17][14] ;
 wire \regs[17][15] ;
 wire \regs[17][16] ;
 wire \regs[17][17] ;
 wire \regs[17][18] ;
 wire \regs[17][19] ;
 wire \regs[17][1] ;
 wire \regs[17][20] ;
 wire \regs[17][21] ;
 wire \regs[17][22] ;
 wire \regs[17][23] ;
 wire \regs[17][24] ;
 wire \regs[17][25] ;
 wire \regs[17][26] ;
 wire \regs[17][27] ;
 wire \regs[17][28] ;
 wire \regs[17][29] ;
 wire \regs[17][2] ;
 wire \regs[17][30] ;
 wire \regs[17][31] ;
 wire \regs[17][3] ;
 wire \regs[17][4] ;
 wire \regs[17][5] ;
 wire \regs[17][6] ;
 wire \regs[17][7] ;
 wire \regs[17][8] ;
 wire \regs[17][9] ;
 wire \regs[18][0] ;
 wire \regs[18][10] ;
 wire \regs[18][11] ;
 wire \regs[18][12] ;
 wire \regs[18][13] ;
 wire \regs[18][14] ;
 wire \regs[18][15] ;
 wire \regs[18][16] ;
 wire \regs[18][17] ;
 wire \regs[18][18] ;
 wire \regs[18][19] ;
 wire \regs[18][1] ;
 wire \regs[18][20] ;
 wire \regs[18][21] ;
 wire \regs[18][22] ;
 wire \regs[18][23] ;
 wire \regs[18][24] ;
 wire \regs[18][25] ;
 wire \regs[18][26] ;
 wire \regs[18][27] ;
 wire \regs[18][28] ;
 wire \regs[18][29] ;
 wire \regs[18][2] ;
 wire \regs[18][30] ;
 wire \regs[18][31] ;
 wire \regs[18][3] ;
 wire \regs[18][4] ;
 wire \regs[18][5] ;
 wire \regs[18][6] ;
 wire \regs[18][7] ;
 wire \regs[18][8] ;
 wire \regs[18][9] ;
 wire \regs[19][0] ;
 wire \regs[19][10] ;
 wire \regs[19][11] ;
 wire \regs[19][12] ;
 wire \regs[19][13] ;
 wire \regs[19][14] ;
 wire \regs[19][15] ;
 wire \regs[19][16] ;
 wire \regs[19][17] ;
 wire \regs[19][18] ;
 wire \regs[19][19] ;
 wire \regs[19][1] ;
 wire \regs[19][20] ;
 wire \regs[19][21] ;
 wire \regs[19][22] ;
 wire \regs[19][23] ;
 wire \regs[19][24] ;
 wire \regs[19][25] ;
 wire \regs[19][26] ;
 wire \regs[19][27] ;
 wire \regs[19][28] ;
 wire \regs[19][29] ;
 wire \regs[19][2] ;
 wire \regs[19][30] ;
 wire \regs[19][31] ;
 wire \regs[19][3] ;
 wire \regs[19][4] ;
 wire \regs[19][5] ;
 wire \regs[19][6] ;
 wire \regs[19][7] ;
 wire \regs[19][8] ;
 wire \regs[19][9] ;
 wire \regs[1][0] ;
 wire \regs[1][10] ;
 wire \regs[1][11] ;
 wire \regs[1][12] ;
 wire \regs[1][13] ;
 wire \regs[1][14] ;
 wire \regs[1][15] ;
 wire \regs[1][16] ;
 wire \regs[1][17] ;
 wire \regs[1][18] ;
 wire \regs[1][19] ;
 wire \regs[1][1] ;
 wire \regs[1][20] ;
 wire \regs[1][21] ;
 wire \regs[1][22] ;
 wire \regs[1][23] ;
 wire \regs[1][24] ;
 wire \regs[1][25] ;
 wire \regs[1][26] ;
 wire \regs[1][27] ;
 wire \regs[1][28] ;
 wire \regs[1][29] ;
 wire \regs[1][2] ;
 wire \regs[1][30] ;
 wire \regs[1][31] ;
 wire \regs[1][3] ;
 wire \regs[1][4] ;
 wire \regs[1][5] ;
 wire \regs[1][6] ;
 wire \regs[1][7] ;
 wire \regs[1][8] ;
 wire \regs[1][9] ;
 wire \regs[20][0] ;
 wire \regs[20][10] ;
 wire \regs[20][11] ;
 wire \regs[20][12] ;
 wire \regs[20][13] ;
 wire \regs[20][14] ;
 wire \regs[20][15] ;
 wire \regs[20][16] ;
 wire \regs[20][17] ;
 wire \regs[20][18] ;
 wire \regs[20][19] ;
 wire \regs[20][1] ;
 wire \regs[20][20] ;
 wire \regs[20][21] ;
 wire \regs[20][22] ;
 wire \regs[20][23] ;
 wire \regs[20][24] ;
 wire \regs[20][25] ;
 wire \regs[20][26] ;
 wire \regs[20][27] ;
 wire \regs[20][28] ;
 wire \regs[20][29] ;
 wire \regs[20][2] ;
 wire \regs[20][30] ;
 wire \regs[20][31] ;
 wire \regs[20][3] ;
 wire \regs[20][4] ;
 wire \regs[20][5] ;
 wire \regs[20][6] ;
 wire \regs[20][7] ;
 wire \regs[20][8] ;
 wire \regs[20][9] ;
 wire \regs[21][0] ;
 wire \regs[21][10] ;
 wire \regs[21][11] ;
 wire \regs[21][12] ;
 wire \regs[21][13] ;
 wire \regs[21][14] ;
 wire \regs[21][15] ;
 wire \regs[21][16] ;
 wire \regs[21][17] ;
 wire \regs[21][18] ;
 wire \regs[21][19] ;
 wire \regs[21][1] ;
 wire \regs[21][20] ;
 wire \regs[21][21] ;
 wire \regs[21][22] ;
 wire \regs[21][23] ;
 wire \regs[21][24] ;
 wire \regs[21][25] ;
 wire \regs[21][26] ;
 wire \regs[21][27] ;
 wire \regs[21][28] ;
 wire \regs[21][29] ;
 wire \regs[21][2] ;
 wire \regs[21][30] ;
 wire \regs[21][31] ;
 wire \regs[21][3] ;
 wire \regs[21][4] ;
 wire \regs[21][5] ;
 wire \regs[21][6] ;
 wire \regs[21][7] ;
 wire \regs[21][8] ;
 wire \regs[21][9] ;
 wire \regs[22][0] ;
 wire \regs[22][10] ;
 wire \regs[22][11] ;
 wire \regs[22][12] ;
 wire \regs[22][13] ;
 wire \regs[22][14] ;
 wire \regs[22][15] ;
 wire \regs[22][16] ;
 wire \regs[22][17] ;
 wire \regs[22][18] ;
 wire \regs[22][19] ;
 wire \regs[22][1] ;
 wire \regs[22][20] ;
 wire \regs[22][21] ;
 wire \regs[22][22] ;
 wire \regs[22][23] ;
 wire \regs[22][24] ;
 wire \regs[22][25] ;
 wire \regs[22][26] ;
 wire \regs[22][27] ;
 wire \regs[22][28] ;
 wire \regs[22][29] ;
 wire \regs[22][2] ;
 wire \regs[22][30] ;
 wire \regs[22][31] ;
 wire \regs[22][3] ;
 wire \regs[22][4] ;
 wire \regs[22][5] ;
 wire \regs[22][6] ;
 wire \regs[22][7] ;
 wire \regs[22][8] ;
 wire \regs[22][9] ;
 wire \regs[23][0] ;
 wire \regs[23][10] ;
 wire \regs[23][11] ;
 wire \regs[23][12] ;
 wire \regs[23][13] ;
 wire \regs[23][14] ;
 wire \regs[23][15] ;
 wire \regs[23][16] ;
 wire \regs[23][17] ;
 wire \regs[23][18] ;
 wire \regs[23][19] ;
 wire \regs[23][1] ;
 wire \regs[23][20] ;
 wire \regs[23][21] ;
 wire \regs[23][22] ;
 wire \regs[23][23] ;
 wire \regs[23][24] ;
 wire \regs[23][25] ;
 wire \regs[23][26] ;
 wire \regs[23][27] ;
 wire \regs[23][28] ;
 wire \regs[23][29] ;
 wire \regs[23][2] ;
 wire \regs[23][30] ;
 wire \regs[23][31] ;
 wire \regs[23][3] ;
 wire \regs[23][4] ;
 wire \regs[23][5] ;
 wire \regs[23][6] ;
 wire \regs[23][7] ;
 wire \regs[23][8] ;
 wire \regs[23][9] ;
 wire \regs[24][0] ;
 wire \regs[24][10] ;
 wire \regs[24][11] ;
 wire \regs[24][12] ;
 wire \regs[24][13] ;
 wire \regs[24][14] ;
 wire \regs[24][15] ;
 wire \regs[24][16] ;
 wire \regs[24][17] ;
 wire \regs[24][18] ;
 wire \regs[24][19] ;
 wire \regs[24][1] ;
 wire \regs[24][20] ;
 wire \regs[24][21] ;
 wire \regs[24][22] ;
 wire \regs[24][23] ;
 wire \regs[24][24] ;
 wire \regs[24][25] ;
 wire \regs[24][26] ;
 wire \regs[24][27] ;
 wire \regs[24][28] ;
 wire \regs[24][29] ;
 wire \regs[24][2] ;
 wire \regs[24][30] ;
 wire \regs[24][31] ;
 wire \regs[24][3] ;
 wire \regs[24][4] ;
 wire \regs[24][5] ;
 wire \regs[24][6] ;
 wire \regs[24][7] ;
 wire \regs[24][8] ;
 wire \regs[24][9] ;
 wire \regs[25][0] ;
 wire \regs[25][10] ;
 wire \regs[25][11] ;
 wire \regs[25][12] ;
 wire \regs[25][13] ;
 wire \regs[25][14] ;
 wire \regs[25][15] ;
 wire \regs[25][16] ;
 wire \regs[25][17] ;
 wire \regs[25][18] ;
 wire \regs[25][19] ;
 wire \regs[25][1] ;
 wire \regs[25][20] ;
 wire \regs[25][21] ;
 wire \regs[25][22] ;
 wire \regs[25][23] ;
 wire \regs[25][24] ;
 wire \regs[25][25] ;
 wire \regs[25][26] ;
 wire \regs[25][27] ;
 wire \regs[25][28] ;
 wire \regs[25][29] ;
 wire \regs[25][2] ;
 wire \regs[25][30] ;
 wire \regs[25][31] ;
 wire \regs[25][3] ;
 wire \regs[25][4] ;
 wire \regs[25][5] ;
 wire \regs[25][6] ;
 wire \regs[25][7] ;
 wire \regs[25][8] ;
 wire \regs[25][9] ;
 wire \regs[26][0] ;
 wire \regs[26][10] ;
 wire \regs[26][11] ;
 wire \regs[26][12] ;
 wire \regs[26][13] ;
 wire \regs[26][14] ;
 wire \regs[26][15] ;
 wire \regs[26][16] ;
 wire \regs[26][17] ;
 wire \regs[26][18] ;
 wire \regs[26][19] ;
 wire \regs[26][1] ;
 wire \regs[26][20] ;
 wire \regs[26][21] ;
 wire \regs[26][22] ;
 wire \regs[26][23] ;
 wire \regs[26][24] ;
 wire \regs[26][25] ;
 wire \regs[26][26] ;
 wire \regs[26][27] ;
 wire \regs[26][28] ;
 wire \regs[26][29] ;
 wire \regs[26][2] ;
 wire \regs[26][30] ;
 wire \regs[26][31] ;
 wire \regs[26][3] ;
 wire \regs[26][4] ;
 wire \regs[26][5] ;
 wire \regs[26][6] ;
 wire \regs[26][7] ;
 wire \regs[26][8] ;
 wire \regs[26][9] ;
 wire \regs[27][0] ;
 wire \regs[27][10] ;
 wire \regs[27][11] ;
 wire \regs[27][12] ;
 wire \regs[27][13] ;
 wire \regs[27][14] ;
 wire \regs[27][15] ;
 wire \regs[27][16] ;
 wire \regs[27][17] ;
 wire \regs[27][18] ;
 wire \regs[27][19] ;
 wire \regs[27][1] ;
 wire \regs[27][20] ;
 wire \regs[27][21] ;
 wire \regs[27][22] ;
 wire \regs[27][23] ;
 wire \regs[27][24] ;
 wire \regs[27][25] ;
 wire \regs[27][26] ;
 wire \regs[27][27] ;
 wire \regs[27][28] ;
 wire \regs[27][29] ;
 wire \regs[27][2] ;
 wire \regs[27][30] ;
 wire \regs[27][31] ;
 wire \regs[27][3] ;
 wire \regs[27][4] ;
 wire \regs[27][5] ;
 wire \regs[27][6] ;
 wire \regs[27][7] ;
 wire \regs[27][8] ;
 wire \regs[27][9] ;
 wire \regs[28][0] ;
 wire \regs[28][10] ;
 wire \regs[28][11] ;
 wire \regs[28][12] ;
 wire \regs[28][13] ;
 wire \regs[28][14] ;
 wire \regs[28][15] ;
 wire \regs[28][16] ;
 wire \regs[28][17] ;
 wire \regs[28][18] ;
 wire \regs[28][19] ;
 wire \regs[28][1] ;
 wire \regs[28][20] ;
 wire \regs[28][21] ;
 wire \regs[28][22] ;
 wire \regs[28][23] ;
 wire \regs[28][24] ;
 wire \regs[28][25] ;
 wire \regs[28][26] ;
 wire \regs[28][27] ;
 wire \regs[28][28] ;
 wire \regs[28][29] ;
 wire \regs[28][2] ;
 wire \regs[28][30] ;
 wire \regs[28][31] ;
 wire \regs[28][3] ;
 wire \regs[28][4] ;
 wire \regs[28][5] ;
 wire \regs[28][6] ;
 wire \regs[28][7] ;
 wire \regs[28][8] ;
 wire \regs[28][9] ;
 wire \regs[29][0] ;
 wire \regs[29][10] ;
 wire \regs[29][11] ;
 wire \regs[29][12] ;
 wire \regs[29][13] ;
 wire \regs[29][14] ;
 wire \regs[29][15] ;
 wire \regs[29][16] ;
 wire \regs[29][17] ;
 wire \regs[29][18] ;
 wire \regs[29][19] ;
 wire \regs[29][1] ;
 wire \regs[29][20] ;
 wire \regs[29][21] ;
 wire \regs[29][22] ;
 wire \regs[29][23] ;
 wire \regs[29][24] ;
 wire \regs[29][25] ;
 wire \regs[29][26] ;
 wire \regs[29][27] ;
 wire \regs[29][28] ;
 wire \regs[29][29] ;
 wire \regs[29][2] ;
 wire \regs[29][30] ;
 wire \regs[29][31] ;
 wire \regs[29][3] ;
 wire \regs[29][4] ;
 wire \regs[29][5] ;
 wire \regs[29][6] ;
 wire \regs[29][7] ;
 wire \regs[29][8] ;
 wire \regs[29][9] ;
 wire \regs[2][0] ;
 wire \regs[2][10] ;
 wire \regs[2][11] ;
 wire \regs[2][12] ;
 wire \regs[2][13] ;
 wire \regs[2][14] ;
 wire \regs[2][15] ;
 wire \regs[2][16] ;
 wire \regs[2][17] ;
 wire \regs[2][18] ;
 wire \regs[2][19] ;
 wire \regs[2][1] ;
 wire \regs[2][20] ;
 wire \regs[2][21] ;
 wire \regs[2][22] ;
 wire \regs[2][23] ;
 wire \regs[2][24] ;
 wire \regs[2][25] ;
 wire \regs[2][26] ;
 wire \regs[2][27] ;
 wire \regs[2][28] ;
 wire \regs[2][29] ;
 wire \regs[2][2] ;
 wire \regs[2][30] ;
 wire \regs[2][31] ;
 wire \regs[2][3] ;
 wire \regs[2][4] ;
 wire \regs[2][5] ;
 wire \regs[2][6] ;
 wire \regs[2][7] ;
 wire \regs[2][8] ;
 wire \regs[2][9] ;
 wire \regs[30][0] ;
 wire \regs[30][10] ;
 wire \regs[30][11] ;
 wire \regs[30][12] ;
 wire \regs[30][13] ;
 wire \regs[30][14] ;
 wire \regs[30][15] ;
 wire \regs[30][16] ;
 wire \regs[30][17] ;
 wire \regs[30][18] ;
 wire \regs[30][19] ;
 wire \regs[30][1] ;
 wire \regs[30][20] ;
 wire \regs[30][21] ;
 wire \regs[30][22] ;
 wire \regs[30][23] ;
 wire \regs[30][24] ;
 wire \regs[30][25] ;
 wire \regs[30][26] ;
 wire \regs[30][27] ;
 wire \regs[30][28] ;
 wire \regs[30][29] ;
 wire \regs[30][2] ;
 wire \regs[30][30] ;
 wire \regs[30][31] ;
 wire \regs[30][3] ;
 wire \regs[30][4] ;
 wire \regs[30][5] ;
 wire \regs[30][6] ;
 wire \regs[30][7] ;
 wire \regs[30][8] ;
 wire \regs[30][9] ;
 wire \regs[31][0] ;
 wire \regs[31][10] ;
 wire \regs[31][11] ;
 wire \regs[31][12] ;
 wire \regs[31][13] ;
 wire \regs[31][14] ;
 wire \regs[31][15] ;
 wire \regs[31][16] ;
 wire \regs[31][17] ;
 wire \regs[31][18] ;
 wire \regs[31][19] ;
 wire \regs[31][1] ;
 wire \regs[31][20] ;
 wire \regs[31][21] ;
 wire \regs[31][22] ;
 wire \regs[31][23] ;
 wire \regs[31][24] ;
 wire \regs[31][25] ;
 wire \regs[31][26] ;
 wire \regs[31][27] ;
 wire \regs[31][28] ;
 wire \regs[31][29] ;
 wire \regs[31][2] ;
 wire \regs[31][30] ;
 wire \regs[31][31] ;
 wire \regs[31][3] ;
 wire \regs[31][4] ;
 wire \regs[31][5] ;
 wire \regs[31][6] ;
 wire \regs[31][7] ;
 wire \regs[31][8] ;
 wire \regs[31][9] ;
 wire \regs[3][0] ;
 wire \regs[3][10] ;
 wire \regs[3][11] ;
 wire \regs[3][12] ;
 wire \regs[3][13] ;
 wire \regs[3][14] ;
 wire \regs[3][15] ;
 wire \regs[3][16] ;
 wire \regs[3][17] ;
 wire \regs[3][18] ;
 wire \regs[3][19] ;
 wire \regs[3][1] ;
 wire \regs[3][20] ;
 wire \regs[3][21] ;
 wire \regs[3][22] ;
 wire \regs[3][23] ;
 wire \regs[3][24] ;
 wire \regs[3][25] ;
 wire \regs[3][26] ;
 wire \regs[3][27] ;
 wire \regs[3][28] ;
 wire \regs[3][29] ;
 wire \regs[3][2] ;
 wire \regs[3][30] ;
 wire \regs[3][31] ;
 wire \regs[3][3] ;
 wire \regs[3][4] ;
 wire \regs[3][5] ;
 wire \regs[3][6] ;
 wire \regs[3][7] ;
 wire \regs[3][8] ;
 wire \regs[3][9] ;
 wire \regs[4][0] ;
 wire \regs[4][10] ;
 wire \regs[4][11] ;
 wire \regs[4][12] ;
 wire \regs[4][13] ;
 wire \regs[4][14] ;
 wire \regs[4][15] ;
 wire \regs[4][16] ;
 wire \regs[4][17] ;
 wire \regs[4][18] ;
 wire \regs[4][19] ;
 wire \regs[4][1] ;
 wire \regs[4][20] ;
 wire \regs[4][21] ;
 wire \regs[4][22] ;
 wire \regs[4][23] ;
 wire \regs[4][24] ;
 wire \regs[4][25] ;
 wire \regs[4][26] ;
 wire \regs[4][27] ;
 wire \regs[4][28] ;
 wire \regs[4][29] ;
 wire \regs[4][2] ;
 wire \regs[4][30] ;
 wire \regs[4][31] ;
 wire \regs[4][3] ;
 wire \regs[4][4] ;
 wire \regs[4][5] ;
 wire \regs[4][6] ;
 wire \regs[4][7] ;
 wire \regs[4][8] ;
 wire \regs[4][9] ;
 wire \regs[5][0] ;
 wire \regs[5][10] ;
 wire \regs[5][11] ;
 wire \regs[5][12] ;
 wire \regs[5][13] ;
 wire \regs[5][14] ;
 wire \regs[5][15] ;
 wire \regs[5][16] ;
 wire \regs[5][17] ;
 wire \regs[5][18] ;
 wire \regs[5][19] ;
 wire \regs[5][1] ;
 wire \regs[5][20] ;
 wire \regs[5][21] ;
 wire \regs[5][22] ;
 wire \regs[5][23] ;
 wire \regs[5][24] ;
 wire \regs[5][25] ;
 wire \regs[5][26] ;
 wire \regs[5][27] ;
 wire \regs[5][28] ;
 wire \regs[5][29] ;
 wire \regs[5][2] ;
 wire \regs[5][30] ;
 wire \regs[5][31] ;
 wire \regs[5][3] ;
 wire \regs[5][4] ;
 wire \regs[5][5] ;
 wire \regs[5][6] ;
 wire \regs[5][7] ;
 wire \regs[5][8] ;
 wire \regs[5][9] ;
 wire \regs[6][0] ;
 wire \regs[6][10] ;
 wire \regs[6][11] ;
 wire \regs[6][12] ;
 wire \regs[6][13] ;
 wire \regs[6][14] ;
 wire \regs[6][15] ;
 wire \regs[6][16] ;
 wire \regs[6][17] ;
 wire \regs[6][18] ;
 wire \regs[6][19] ;
 wire \regs[6][1] ;
 wire \regs[6][20] ;
 wire \regs[6][21] ;
 wire \regs[6][22] ;
 wire \regs[6][23] ;
 wire \regs[6][24] ;
 wire \regs[6][25] ;
 wire \regs[6][26] ;
 wire \regs[6][27] ;
 wire \regs[6][28] ;
 wire \regs[6][29] ;
 wire \regs[6][2] ;
 wire \regs[6][30] ;
 wire \regs[6][31] ;
 wire \regs[6][3] ;
 wire \regs[6][4] ;
 wire \regs[6][5] ;
 wire \regs[6][6] ;
 wire \regs[6][7] ;
 wire \regs[6][8] ;
 wire \regs[6][9] ;
 wire \regs[7][0] ;
 wire \regs[7][10] ;
 wire \regs[7][11] ;
 wire \regs[7][12] ;
 wire \regs[7][13] ;
 wire \regs[7][14] ;
 wire \regs[7][15] ;
 wire \regs[7][16] ;
 wire \regs[7][17] ;
 wire \regs[7][18] ;
 wire \regs[7][19] ;
 wire \regs[7][1] ;
 wire \regs[7][20] ;
 wire \regs[7][21] ;
 wire \regs[7][22] ;
 wire \regs[7][23] ;
 wire \regs[7][24] ;
 wire \regs[7][25] ;
 wire \regs[7][26] ;
 wire \regs[7][27] ;
 wire \regs[7][28] ;
 wire \regs[7][29] ;
 wire \regs[7][2] ;
 wire \regs[7][30] ;
 wire \regs[7][31] ;
 wire \regs[7][3] ;
 wire \regs[7][4] ;
 wire \regs[7][5] ;
 wire \regs[7][6] ;
 wire \regs[7][7] ;
 wire \regs[7][8] ;
 wire \regs[7][9] ;
 wire \regs[8][0] ;
 wire \regs[8][10] ;
 wire \regs[8][11] ;
 wire \regs[8][12] ;
 wire \regs[8][13] ;
 wire \regs[8][14] ;
 wire \regs[8][15] ;
 wire \regs[8][16] ;
 wire \regs[8][17] ;
 wire \regs[8][18] ;
 wire \regs[8][19] ;
 wire \regs[8][1] ;
 wire \regs[8][20] ;
 wire \regs[8][21] ;
 wire \regs[8][22] ;
 wire \regs[8][23] ;
 wire \regs[8][24] ;
 wire \regs[8][25] ;
 wire \regs[8][26] ;
 wire \regs[8][27] ;
 wire \regs[8][28] ;
 wire \regs[8][29] ;
 wire \regs[8][2] ;
 wire \regs[8][30] ;
 wire \regs[8][31] ;
 wire \regs[8][3] ;
 wire \regs[8][4] ;
 wire \regs[8][5] ;
 wire \regs[8][6] ;
 wire \regs[8][7] ;
 wire \regs[8][8] ;
 wire \regs[8][9] ;
 wire \regs[9][0] ;
 wire \regs[9][10] ;
 wire \regs[9][11] ;
 wire \regs[9][12] ;
 wire \regs[9][13] ;
 wire \regs[9][14] ;
 wire \regs[9][15] ;
 wire \regs[9][16] ;
 wire \regs[9][17] ;
 wire \regs[9][18] ;
 wire \regs[9][19] ;
 wire \regs[9][1] ;
 wire \regs[9][20] ;
 wire \regs[9][21] ;
 wire \regs[9][22] ;
 wire \regs[9][23] ;
 wire \regs[9][24] ;
 wire \regs[9][25] ;
 wire \regs[9][26] ;
 wire \regs[9][27] ;
 wire \regs[9][28] ;
 wire \regs[9][29] ;
 wire \regs[9][2] ;
 wire \regs[9][30] ;
 wire \regs[9][31] ;
 wire \regs[9][3] ;
 wire \regs[9][4] ;
 wire \regs[9][5] ;
 wire \regs[9][6] ;
 wire \regs[9][7] ;
 wire \regs[9][8] ;
 wire \regs[9][9] ;
 wire \rs2_content[0] ;
 wire \rs2_content[10] ;
 wire \rs2_content[11] ;
 wire \rs2_content[12] ;
 wire \rs2_content[13] ;
 wire \rs2_content[14] ;
 wire \rs2_content[15] ;
 wire \rs2_content[16] ;
 wire \rs2_content[17] ;
 wire \rs2_content[18] ;
 wire \rs2_content[19] ;
 wire \rs2_content[1] ;
 wire \rs2_content[20] ;
 wire \rs2_content[21] ;
 wire \rs2_content[22] ;
 wire \rs2_content[23] ;
 wire \rs2_content[24] ;
 wire \rs2_content[25] ;
 wire \rs2_content[26] ;
 wire \rs2_content[27] ;
 wire \rs2_content[28] ;
 wire \rs2_content[29] ;
 wire \rs2_content[2] ;
 wire \rs2_content[30] ;
 wire \rs2_content[31] ;
 wire \rs2_content[3] ;
 wire \rs2_content[4] ;
 wire \rs2_content[5] ;
 wire \rs2_content[6] ;
 wire \rs2_content[7] ;
 wire \rs2_content[8] ;
 wire \rs2_content[9] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_59_clk;
 wire clknet_leaf_60_clk;
 wire clknet_leaf_61_clk;
 wire clknet_leaf_62_clk;
 wire clknet_leaf_63_clk;
 wire clknet_leaf_64_clk;
 wire clknet_leaf_65_clk;
 wire clknet_leaf_66_clk;
 wire clknet_leaf_67_clk;
 wire clknet_leaf_68_clk;
 wire clknet_leaf_69_clk;
 wire clknet_leaf_70_clk;
 wire clknet_leaf_71_clk;
 wire clknet_leaf_72_clk;
 wire clknet_leaf_73_clk;
 wire clknet_leaf_74_clk;
 wire clknet_leaf_75_clk;
 wire clknet_leaf_76_clk;
 wire clknet_leaf_77_clk;
 wire clknet_leaf_78_clk;
 wire clknet_leaf_79_clk;
 wire clknet_leaf_80_clk;
 wire clknet_leaf_81_clk;
 wire clknet_leaf_82_clk;
 wire clknet_leaf_83_clk;
 wire clknet_leaf_84_clk;
 wire clknet_leaf_85_clk;
 wire clknet_leaf_86_clk;
 wire clknet_leaf_87_clk;
 wire clknet_leaf_88_clk;
 wire clknet_leaf_89_clk;
 wire clknet_leaf_90_clk;
 wire clknet_leaf_91_clk;
 wire clknet_leaf_92_clk;
 wire clknet_leaf_93_clk;
 wire clknet_leaf_94_clk;
 wire clknet_leaf_95_clk;
 wire clknet_leaf_96_clk;
 wire clknet_leaf_97_clk;
 wire clknet_leaf_98_clk;
 wire clknet_leaf_99_clk;
 wire clknet_leaf_100_clk;
 wire clknet_leaf_101_clk;
 wire clknet_leaf_102_clk;
 wire clknet_leaf_103_clk;
 wire clknet_leaf_104_clk;
 wire clknet_leaf_105_clk;
 wire clknet_leaf_106_clk;
 wire clknet_leaf_107_clk;
 wire clknet_leaf_108_clk;
 wire clknet_leaf_109_clk;
 wire clknet_leaf_110_clk;
 wire clknet_leaf_111_clk;
 wire clknet_leaf_112_clk;
 wire clknet_leaf_113_clk;
 wire clknet_leaf_114_clk;
 wire clknet_leaf_115_clk;
 wire clknet_leaf_116_clk;
 wire clknet_leaf_117_clk;
 wire clknet_leaf_118_clk;
 wire clknet_leaf_119_clk;
 wire clknet_leaf_120_clk;
 wire clknet_leaf_121_clk;
 wire clknet_leaf_122_clk;
 wire clknet_leaf_123_clk;
 wire clknet_leaf_124_clk;
 wire clknet_leaf_125_clk;
 wire clknet_leaf_126_clk;
 wire clknet_leaf_127_clk;
 wire clknet_leaf_128_clk;
 wire clknet_leaf_129_clk;
 wire clknet_leaf_130_clk;
 wire clknet_leaf_131_clk;
 wire clknet_leaf_132_clk;
 wire clknet_leaf_133_clk;
 wire clknet_leaf_134_clk;
 wire clknet_leaf_135_clk;
 wire clknet_0_clk;
 wire clknet_1_0_0_clk;
 wire clknet_1_1_0_clk;
 wire clknet_2_0_0_clk;
 wire clknet_2_1_0_clk;
 wire clknet_2_2_0_clk;
 wire clknet_2_3_0_clk;
 wire clknet_3_0_0_clk;
 wire clknet_3_1_0_clk;
 wire clknet_3_2_0_clk;
 wire clknet_3_3_0_clk;
 wire clknet_3_4_0_clk;
 wire clknet_3_5_0_clk;
 wire clknet_3_6_0_clk;
 wire clknet_3_7_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_opt_1_0_clk;
 wire clknet_opt_2_0_clk;
 wire clknet_opt_3_0_clk;

 sky130_fd_sc_hd__inv_2 _07032_ (.A(\core_state[1] ),
    .Y(_01526_));
 sky130_fd_sc_hd__clkbuf_4 _07033_ (.A(_01526_),
    .X(_01527_));
 sky130_fd_sc_hd__clkbuf_4 _07034_ (.A(_01527_),
    .X(_01528_));
 sky130_fd_sc_hd__buf_4 _07035_ (.A(_01528_),
    .X(_01529_));
 sky130_fd_sc_hd__buf_2 _07036_ (.A(\instr[4] ),
    .X(_01530_));
 sky130_fd_sc_hd__and3b_2 _07037_ (.A_N(_01530_),
    .B(\instr[5] ),
    .C(\instr[6] ),
    .X(_01531_));
 sky130_fd_sc_hd__and4_4 _07038_ (.A(\instr[2] ),
    .B(\instr[1] ),
    .C(\instr[0] ),
    .D(_01531_),
    .X(_01532_));
 sky130_fd_sc_hd__and2_1 _07039_ (.A(\instr[3] ),
    .B(_01532_),
    .X(_01533_));
 sky130_fd_sc_hd__buf_4 _07040_ (.A(_01533_),
    .X(_01534_));
 sky130_fd_sc_hd__buf_6 _07041_ (.A(\B_type_imm[12] ),
    .X(_01535_));
 sky130_fd_sc_hd__buf_4 _07042_ (.A(_01535_),
    .X(_01536_));
 sky130_fd_sc_hd__buf_2 _07043_ (.A(_01536_),
    .X(_01537_));
 sky130_fd_sc_hd__clkbuf_4 _07044_ (.A(_01537_),
    .X(_01538_));
 sky130_fd_sc_hd__clkbuf_4 _07045_ (.A(_01538_),
    .X(_01539_));
 sky130_fd_sc_hd__buf_4 _07046_ (.A(_01539_),
    .X(_01540_));
 sky130_fd_sc_hd__xor2_1 _07047_ (.A(\PC[23] ),
    .B(_01540_),
    .X(_01541_));
 sky130_fd_sc_hd__or2_1 _07048_ (.A(\PC[22] ),
    .B(_01538_),
    .X(_01542_));
 sky130_fd_sc_hd__nand2_1 _07049_ (.A(\PC[21] ),
    .B(_01538_),
    .Y(_01543_));
 sky130_fd_sc_hd__or2_1 _07050_ (.A(\PC[21] ),
    .B(_01538_),
    .X(_01544_));
 sky130_fd_sc_hd__nand2_1 _07051_ (.A(_01543_),
    .B(_01544_),
    .Y(_01545_));
 sky130_fd_sc_hd__clkbuf_4 _07052_ (.A(\PC[20] ),
    .X(_01546_));
 sky130_fd_sc_hd__nand2_1 _07053_ (.A(_01546_),
    .B(_01537_),
    .Y(_01547_));
 sky130_fd_sc_hd__nand2_1 _07054_ (.A(\PC[19] ),
    .B(\J_type_imm[19] ),
    .Y(_01548_));
 sky130_fd_sc_hd__and2_1 _07055_ (.A(\PC[18] ),
    .B(\J_type_imm[18] ),
    .X(_01549_));
 sky130_fd_sc_hd__or2_1 _07056_ (.A(\PC[18] ),
    .B(\J_type_imm[18] ),
    .X(_01550_));
 sky130_fd_sc_hd__and2b_1 _07057_ (.A_N(_01549_),
    .B(_01550_),
    .X(_01551_));
 sky130_fd_sc_hd__and2_1 _07058_ (.A(\PC[17] ),
    .B(\J_type_imm[17] ),
    .X(_01552_));
 sky130_fd_sc_hd__nor2_1 _07059_ (.A(\PC[17] ),
    .B(\J_type_imm[17] ),
    .Y(_01553_));
 sky130_fd_sc_hd__or2_1 _07060_ (.A(_01552_),
    .B(_01553_),
    .X(_01554_));
 sky130_fd_sc_hd__and2_1 _07061_ (.A(\PC[16] ),
    .B(\J_type_imm[16] ),
    .X(_01555_));
 sky130_fd_sc_hd__nor2_1 _07062_ (.A(\PC[16] ),
    .B(\J_type_imm[16] ),
    .Y(_01556_));
 sky130_fd_sc_hd__nor2_1 _07063_ (.A(_01555_),
    .B(_01556_),
    .Y(_01557_));
 sky130_fd_sc_hd__clkbuf_4 _07064_ (.A(\PC[12] ),
    .X(_01558_));
 sky130_fd_sc_hd__and2_1 _07065_ (.A(_01558_),
    .B(\J_type_imm[12] ),
    .X(_01559_));
 sky130_fd_sc_hd__xor2_1 _07066_ (.A(\PC[13] ),
    .B(\J_type_imm[13] ),
    .X(_01560_));
 sky130_fd_sc_hd__and2_1 _07067_ (.A(_01559_),
    .B(_01560_),
    .X(_01561_));
 sky130_fd_sc_hd__inv_2 _07068_ (.A(_01561_),
    .Y(_01562_));
 sky130_fd_sc_hd__nor2_1 _07069_ (.A(_01558_),
    .B(\J_type_imm[12] ),
    .Y(_01563_));
 sky130_fd_sc_hd__clkbuf_4 _07070_ (.A(\I_type_imm[0] ),
    .X(_01564_));
 sky130_fd_sc_hd__nor2_1 _07071_ (.A(\PC[11] ),
    .B(_01564_),
    .Y(_01565_));
 sky130_fd_sc_hd__and2_1 _07072_ (.A(\PC[9] ),
    .B(\B_type_imm[9] ),
    .X(_01566_));
 sky130_fd_sc_hd__clkbuf_4 _07073_ (.A(\B_type_imm[9] ),
    .X(_01567_));
 sky130_fd_sc_hd__nor2_1 _07074_ (.A(\PC[9] ),
    .B(_01567_),
    .Y(_01568_));
 sky130_fd_sc_hd__or2_1 _07075_ (.A(_01566_),
    .B(_01568_),
    .X(_01569_));
 sky130_fd_sc_hd__clkbuf_2 _07076_ (.A(_01569_),
    .X(_01570_));
 sky130_fd_sc_hd__or2_1 _07077_ (.A(\PC[8] ),
    .B(\B_type_imm[8] ),
    .X(_01571_));
 sky130_fd_sc_hd__nand2_2 _07078_ (.A(\PC[8] ),
    .B(\B_type_imm[8] ),
    .Y(_01572_));
 sky130_fd_sc_hd__nand2_2 _07079_ (.A(_01571_),
    .B(_01572_),
    .Y(_01573_));
 sky130_fd_sc_hd__nor2_1 _07080_ (.A(\PC[7] ),
    .B(\B_type_imm[7] ),
    .Y(_01574_));
 sky130_fd_sc_hd__and2_1 _07081_ (.A(\PC[7] ),
    .B(\B_type_imm[7] ),
    .X(_01575_));
 sky130_fd_sc_hd__or2_1 _07082_ (.A(_01574_),
    .B(_01575_),
    .X(_01576_));
 sky130_fd_sc_hd__buf_2 _07083_ (.A(_01576_),
    .X(_01577_));
 sky130_fd_sc_hd__nor2_1 _07084_ (.A(_01573_),
    .B(_01577_),
    .Y(_01578_));
 sky130_fd_sc_hd__or2_1 _07085_ (.A(\PC[4] ),
    .B(\I_type_imm[4] ),
    .X(_01579_));
 sky130_fd_sc_hd__nor2_1 _07086_ (.A(\PC[3] ),
    .B(\I_type_imm[3] ),
    .Y(_01580_));
 sky130_fd_sc_hd__inv_2 _07087_ (.A(_01580_),
    .Y(_01581_));
 sky130_fd_sc_hd__xor2_1 _07088_ (.A(\PC[2] ),
    .B(\I_type_imm[2] ),
    .X(_01582_));
 sky130_fd_sc_hd__and2_1 _07089_ (.A(\I_type_imm[1] ),
    .B(\PC[1] ),
    .X(_01583_));
 sky130_fd_sc_hd__and2_1 _07090_ (.A(\PC[3] ),
    .B(\I_type_imm[3] ),
    .X(_01584_));
 sky130_fd_sc_hd__buf_2 _07091_ (.A(\PC[2] ),
    .X(_01585_));
 sky130_fd_sc_hd__and2_1 _07092_ (.A(_01585_),
    .B(\I_type_imm[2] ),
    .X(_01586_));
 sky130_fd_sc_hd__a211o_1 _07093_ (.A1(_01582_),
    .A2(_01583_),
    .B1(_01584_),
    .C1(_01586_),
    .X(_01587_));
 sky130_fd_sc_hd__and2_1 _07094_ (.A(\PC[4] ),
    .B(\I_type_imm[4] ),
    .X(_01588_));
 sky130_fd_sc_hd__a31o_1 _07095_ (.A1(_01579_),
    .A2(_01581_),
    .A3(_01587_),
    .B1(_01588_),
    .X(_01589_));
 sky130_fd_sc_hd__nand2_1 _07096_ (.A(\PC[5] ),
    .B(\B_type_imm[5] ),
    .Y(_01590_));
 sky130_fd_sc_hd__clkbuf_4 _07097_ (.A(\PC[6] ),
    .X(_01591_));
 sky130_fd_sc_hd__xor2_2 _07098_ (.A(_01591_),
    .B(\B_type_imm[6] ),
    .X(_01592_));
 sky130_fd_sc_hd__or2_1 _07099_ (.A(\PC[5] ),
    .B(\B_type_imm[5] ),
    .X(_01593_));
 sky130_fd_sc_hd__and3_1 _07100_ (.A(_01590_),
    .B(_01592_),
    .C(_01593_),
    .X(_01594_));
 sky130_fd_sc_hd__clkbuf_4 _07101_ (.A(\B_type_imm[6] ),
    .X(_01595_));
 sky130_fd_sc_hd__o211a_1 _07102_ (.A1(_01591_),
    .A2(_01595_),
    .B1(\B_type_imm[5] ),
    .C1(\PC[5] ),
    .X(_01596_));
 sky130_fd_sc_hd__a21oi_4 _07103_ (.A1(_01591_),
    .A2(_01595_),
    .B1(_01596_),
    .Y(_01597_));
 sky130_fd_sc_hd__nand3_1 _07104_ (.A(\PC[7] ),
    .B(\B_type_imm[7] ),
    .C(_01571_),
    .Y(_01598_));
 sky130_fd_sc_hd__o311ai_4 _07105_ (.A1(_01597_),
    .A2(_01573_),
    .A3(_01577_),
    .B1(_01572_),
    .C1(_01598_),
    .Y(_01599_));
 sky130_fd_sc_hd__a31oi_4 _07106_ (.A1(_01578_),
    .A2(_01589_),
    .A3(_01594_),
    .B1(_01599_),
    .Y(_01600_));
 sky130_fd_sc_hd__and2_1 _07107_ (.A(\PC[10] ),
    .B(\barrel_shifter_right.arith ),
    .X(_01601_));
 sky130_fd_sc_hd__clkbuf_4 _07108_ (.A(\barrel_shifter_right.arith ),
    .X(_01602_));
 sky130_fd_sc_hd__nor2_1 _07109_ (.A(\PC[10] ),
    .B(_01602_),
    .Y(_01603_));
 sky130_fd_sc_hd__nor2_1 _07110_ (.A(_01601_),
    .B(_01603_),
    .Y(_01604_));
 sky130_fd_sc_hd__inv_2 _07111_ (.A(_01604_),
    .Y(_01605_));
 sky130_fd_sc_hd__o21ba_1 _07112_ (.A1(_01601_),
    .A2(_01566_),
    .B1_N(_01603_),
    .X(_01606_));
 sky130_fd_sc_hd__inv_2 _07113_ (.A(_01606_),
    .Y(_01607_));
 sky130_fd_sc_hd__o31a_1 _07114_ (.A1(_01570_),
    .A2(_01600_),
    .A3(_01605_),
    .B1(_01607_),
    .X(_01608_));
 sky130_fd_sc_hd__and2_1 _07115_ (.A(\PC[11] ),
    .B(\I_type_imm[0] ),
    .X(_01609_));
 sky130_fd_sc_hd__o21ba_1 _07116_ (.A1(_01565_),
    .A2(_01608_),
    .B1_N(_01609_),
    .X(_01610_));
 sky130_fd_sc_hd__or3b_2 _07117_ (.A(_01563_),
    .B(_01610_),
    .C_N(_01560_),
    .X(_01611_));
 sky130_fd_sc_hd__and2_1 _07118_ (.A(\PC[14] ),
    .B(\J_type_imm[14] ),
    .X(_01612_));
 sky130_fd_sc_hd__nor2_1 _07119_ (.A(\PC[14] ),
    .B(\J_type_imm[14] ),
    .Y(_01613_));
 sky130_fd_sc_hd__or2_1 _07120_ (.A(_01612_),
    .B(_01613_),
    .X(_01614_));
 sky130_fd_sc_hd__buf_2 _07121_ (.A(\PC[15] ),
    .X(_01615_));
 sky130_fd_sc_hd__nand2_1 _07122_ (.A(_01615_),
    .B(\J_type_imm[15] ),
    .Y(_01616_));
 sky130_fd_sc_hd__or2_1 _07123_ (.A(_01615_),
    .B(\J_type_imm[15] ),
    .X(_01617_));
 sky130_fd_sc_hd__nand2_1 _07124_ (.A(_01616_),
    .B(_01617_),
    .Y(_01618_));
 sky130_fd_sc_hd__a211oi_1 _07125_ (.A1(_01562_),
    .A2(_01611_),
    .B1(_01614_),
    .C1(_01618_),
    .Y(_01619_));
 sky130_fd_sc_hd__nor2_1 _07126_ (.A(\PC[15] ),
    .B(\J_type_imm[15] ),
    .Y(_01620_));
 sky130_fd_sc_hd__and2_1 _07127_ (.A(\PC[13] ),
    .B(\J_type_imm[13] ),
    .X(_01621_));
 sky130_fd_sc_hd__a211oi_2 _07128_ (.A1(_01559_),
    .A2(_01560_),
    .B1(_01612_),
    .C1(_01621_),
    .Y(_01622_));
 sky130_fd_sc_hd__o31a_1 _07129_ (.A1(_01613_),
    .A2(_01620_),
    .A3(_01622_),
    .B1(_01616_),
    .X(_01623_));
 sky130_fd_sc_hd__o21bai_2 _07130_ (.A1(_01556_),
    .A2(_01623_),
    .B1_N(_01555_),
    .Y(_01624_));
 sky130_fd_sc_hd__a21oi_1 _07131_ (.A1(_01557_),
    .A2(_01619_),
    .B1(_01624_),
    .Y(_01625_));
 sky130_fd_sc_hd__or2_1 _07132_ (.A(_01554_),
    .B(_01625_),
    .X(_01626_));
 sky130_fd_sc_hd__or2b_1 _07133_ (.A(_01552_),
    .B_N(_01626_),
    .X(_01627_));
 sky130_fd_sc_hd__and2_1 _07134_ (.A(_01551_),
    .B(_01627_),
    .X(_01628_));
 sky130_fd_sc_hd__or2_1 _07135_ (.A(\PC[19] ),
    .B(\J_type_imm[19] ),
    .X(_01629_));
 sky130_fd_sc_hd__nand2_1 _07136_ (.A(_01548_),
    .B(_01629_),
    .Y(_01630_));
 sky130_fd_sc_hd__o21bai_1 _07137_ (.A1(_01549_),
    .A2(_01628_),
    .B1_N(_01630_),
    .Y(_01631_));
 sky130_fd_sc_hd__nor2_1 _07138_ (.A(_01546_),
    .B(_01537_),
    .Y(_01632_));
 sky130_fd_sc_hd__a31o_1 _07139_ (.A1(_01547_),
    .A2(_01548_),
    .A3(_01631_),
    .B1(_01632_),
    .X(_01633_));
 sky130_fd_sc_hd__o21ai_1 _07140_ (.A1(_01545_),
    .A2(_01633_),
    .B1(_01543_),
    .Y(_01634_));
 sky130_fd_sc_hd__and2_1 _07141_ (.A(\PC[22] ),
    .B(_01539_),
    .X(_01635_));
 sky130_fd_sc_hd__a21oi_1 _07142_ (.A1(_01542_),
    .A2(_01634_),
    .B1(_01635_),
    .Y(_01636_));
 sky130_fd_sc_hd__xnor2_1 _07143_ (.A(_01541_),
    .B(_01636_),
    .Y(_01637_));
 sky130_fd_sc_hd__or2b_1 _07144_ (.A(_01632_),
    .B_N(_01547_),
    .X(_01638_));
 sky130_fd_sc_hd__inv_2 _07145_ (.A(_01638_),
    .Y(_01639_));
 sky130_fd_sc_hd__xnor2_1 _07146_ (.A(\PC[18] ),
    .B(_01538_),
    .Y(_01640_));
 sky130_fd_sc_hd__xnor2_1 _07147_ (.A(\PC[14] ),
    .B(_01536_),
    .Y(_01641_));
 sky130_fd_sc_hd__buf_4 _07148_ (.A(\B_type_imm[11] ),
    .X(_01642_));
 sky130_fd_sc_hd__or2_1 _07149_ (.A(\PC[11] ),
    .B(_01642_),
    .X(_01643_));
 sky130_fd_sc_hd__inv_2 _07150_ (.A(_01594_),
    .Y(_01644_));
 sky130_fd_sc_hd__nor2_1 _07151_ (.A(\PC[4] ),
    .B(\B_type_imm[4] ),
    .Y(_01645_));
 sky130_fd_sc_hd__nor2_1 _07152_ (.A(\PC[3] ),
    .B(\B_type_imm[3] ),
    .Y(_01646_));
 sky130_fd_sc_hd__nor2_1 _07153_ (.A(_01585_),
    .B(\B_type_imm[2] ),
    .Y(_01647_));
 sky130_fd_sc_hd__clkbuf_8 _07154_ (.A(\B_type_imm[1] ),
    .X(_01648_));
 sky130_fd_sc_hd__nand2_1 _07155_ (.A(_01648_),
    .B(\PC[1] ),
    .Y(_01649_));
 sky130_fd_sc_hd__nand2_1 _07156_ (.A(\PC[3] ),
    .B(\B_type_imm[3] ),
    .Y(_01650_));
 sky130_fd_sc_hd__nand2_1 _07157_ (.A(_01585_),
    .B(\B_type_imm[2] ),
    .Y(_01651_));
 sky130_fd_sc_hd__o211a_1 _07158_ (.A1(_01647_),
    .A2(_01649_),
    .B1(_01650_),
    .C1(_01651_),
    .X(_01652_));
 sky130_fd_sc_hd__nand2_1 _07159_ (.A(\PC[4] ),
    .B(\B_type_imm[4] ),
    .Y(_01653_));
 sky130_fd_sc_hd__o31a_2 _07160_ (.A1(_01645_),
    .A2(_01646_),
    .A3(_01652_),
    .B1(_01653_),
    .X(_01654_));
 sky130_fd_sc_hd__o311a_1 _07161_ (.A1(_01597_),
    .A2(_01573_),
    .A3(_01577_),
    .B1(_01572_),
    .C1(_01598_),
    .X(_01655_));
 sky130_fd_sc_hd__o41a_2 _07162_ (.A1(_01573_),
    .A2(_01577_),
    .A3(_01644_),
    .A4(_01654_),
    .B1(_01655_),
    .X(_01656_));
 sky130_fd_sc_hd__o31ai_2 _07163_ (.A1(_01570_),
    .A2(_01605_),
    .A3(_01656_),
    .B1(_01607_),
    .Y(_01657_));
 sky130_fd_sc_hd__nand2_1 _07164_ (.A(\PC[11] ),
    .B(\B_type_imm[11] ),
    .Y(_01658_));
 sky130_fd_sc_hd__inv_2 _07165_ (.A(_01658_),
    .Y(_01659_));
 sky130_fd_sc_hd__a221o_1 _07166_ (.A1(_01558_),
    .A2(_01535_),
    .B1(_01643_),
    .B2(_01657_),
    .C1(_01659_),
    .X(_01660_));
 sky130_fd_sc_hd__o21a_1 _07167_ (.A1(_01558_),
    .A2(_01535_),
    .B1(_01660_),
    .X(_01661_));
 sky130_fd_sc_hd__nand2_1 _07168_ (.A(\PC[13] ),
    .B(_01535_),
    .Y(_01662_));
 sky130_fd_sc_hd__or2_1 _07169_ (.A(\PC[13] ),
    .B(_01535_),
    .X(_01663_));
 sky130_fd_sc_hd__and2_1 _07170_ (.A(_01662_),
    .B(_01663_),
    .X(_01664_));
 sky130_fd_sc_hd__nand2_1 _07171_ (.A(_01661_),
    .B(_01664_),
    .Y(_01665_));
 sky130_fd_sc_hd__or2_1 _07172_ (.A(_01641_),
    .B(_01665_),
    .X(_01666_));
 sky130_fd_sc_hd__xnor2_1 _07173_ (.A(\PC[16] ),
    .B(_01536_),
    .Y(_01667_));
 sky130_fd_sc_hd__xnor2_1 _07174_ (.A(_01615_),
    .B(_01536_),
    .Y(_01668_));
 sky130_fd_sc_hd__or3_1 _07175_ (.A(_01666_),
    .B(_01667_),
    .C(_01668_),
    .X(_01669_));
 sky130_fd_sc_hd__o21ai_1 _07176_ (.A1(\PC[14] ),
    .A2(\PC[13] ),
    .B1(_01537_),
    .Y(_01670_));
 sky130_fd_sc_hd__o21ai_1 _07177_ (.A1(\PC[16] ),
    .A2(_01615_),
    .B1(_01537_),
    .Y(_01671_));
 sky130_fd_sc_hd__nor2_1 _07178_ (.A(\PC[17] ),
    .B(_01537_),
    .Y(_01672_));
 sky130_fd_sc_hd__and2_1 _07179_ (.A(\PC[17] ),
    .B(_01537_),
    .X(_01673_));
 sky130_fd_sc_hd__a311o_1 _07180_ (.A1(_01669_),
    .A2(_01670_),
    .A3(_01671_),
    .B1(_01672_),
    .C1(_01673_),
    .X(_01674_));
 sky130_fd_sc_hd__nor2_1 _07181_ (.A(_01640_),
    .B(_01674_),
    .Y(_01675_));
 sky130_fd_sc_hd__nand2_1 _07182_ (.A(\PC[19] ),
    .B(_01538_),
    .Y(_01676_));
 sky130_fd_sc_hd__or2_1 _07183_ (.A(\PC[19] ),
    .B(_01537_),
    .X(_01677_));
 sky130_fd_sc_hd__and2_1 _07184_ (.A(_01676_),
    .B(_01677_),
    .X(_01678_));
 sky130_fd_sc_hd__o21a_1 _07185_ (.A1(\PC[18] ),
    .A2(\PC[17] ),
    .B1(_01538_),
    .X(_01679_));
 sky130_fd_sc_hd__nand3b_1 _07186_ (.A_N(_01679_),
    .B(_01676_),
    .C(_01547_),
    .Y(_01680_));
 sky130_fd_sc_hd__a31oi_2 _07187_ (.A1(_01639_),
    .A2(_01675_),
    .A3(_01678_),
    .B1(_01680_),
    .Y(_01681_));
 sky130_fd_sc_hd__o21ai_1 _07188_ (.A1(_01545_),
    .A2(_01681_),
    .B1(_01543_),
    .Y(_01682_));
 sky130_fd_sc_hd__a21oi_1 _07189_ (.A1(_01542_),
    .A2(_01682_),
    .B1(_01635_),
    .Y(_01683_));
 sky130_fd_sc_hd__or2_1 _07190_ (.A(_01541_),
    .B(_01683_),
    .X(_01684_));
 sky130_fd_sc_hd__clkbuf_4 _07191_ (.A(\J_type_imm[14] ),
    .X(_01685_));
 sky130_fd_sc_hd__clkbuf_4 _07192_ (.A(_01685_),
    .X(_01686_));
 sky130_fd_sc_hd__buf_4 _07193_ (.A(_01686_),
    .X(_01687_));
 sky130_fd_sc_hd__inv_6 _07194_ (.A(_01687_),
    .Y(_01688_));
 sky130_fd_sc_hd__buf_6 _07195_ (.A(\J_type_imm[13] ),
    .X(_01689_));
 sky130_fd_sc_hd__and2_2 _07196_ (.A(_01688_),
    .B(_01689_),
    .X(_01690_));
 sky130_fd_sc_hd__and2b_1 _07197_ (.A_N(\leorv32_alu.input1[31] ),
    .B(\rs2_content[31] ),
    .X(_01691_));
 sky130_fd_sc_hd__inv_2 _07198_ (.A(\rs2_content[30] ),
    .Y(_01692_));
 sky130_fd_sc_hd__inv_2 _07199_ (.A(\rs2_content[29] ),
    .Y(_01693_));
 sky130_fd_sc_hd__inv_2 _07200_ (.A(\leorv32_alu.input1[30] ),
    .Y(_01694_));
 sky130_fd_sc_hd__and2b_1 _07201_ (.A_N(\rs2_content[31] ),
    .B(\leorv32_alu.input1[31] ),
    .X(_01695_));
 sky130_fd_sc_hd__a211o_1 _07202_ (.A1(_01694_),
    .A2(\rs2_content[30] ),
    .B1(_01691_),
    .C1(_01695_),
    .X(_01696_));
 sky130_fd_sc_hd__a221o_1 _07203_ (.A1(\leorv32_alu.input1[30] ),
    .A2(_01692_),
    .B1(_01693_),
    .B2(\leorv32_alu.input1[29] ),
    .C1(_01696_),
    .X(_01697_));
 sky130_fd_sc_hd__inv_2 _07204_ (.A(\rs2_content[28] ),
    .Y(_01698_));
 sky130_fd_sc_hd__o22a_1 _07205_ (.A1(\leorv32_alu.input1[29] ),
    .A2(_01693_),
    .B1(_01698_),
    .B2(\leorv32_alu.input1[28] ),
    .X(_01699_));
 sky130_fd_sc_hd__inv_2 _07206_ (.A(\leorv32_alu.input1[27] ),
    .Y(_01700_));
 sky130_fd_sc_hd__nor2_1 _07207_ (.A(_01700_),
    .B(\rs2_content[27] ),
    .Y(_01701_));
 sky130_fd_sc_hd__inv_2 _07208_ (.A(\leorv32_alu.input1[25] ),
    .Y(_01702_));
 sky130_fd_sc_hd__inv_2 _07209_ (.A(\leorv32_alu.input1[24] ),
    .Y(_01703_));
 sky130_fd_sc_hd__a22o_1 _07210_ (.A1(_01702_),
    .A2(\rs2_content[25] ),
    .B1(\rs2_content[24] ),
    .B2(_01703_),
    .X(_01704_));
 sky130_fd_sc_hd__inv_2 _07211_ (.A(\leorv32_alu.input1[26] ),
    .Y(_01705_));
 sky130_fd_sc_hd__o22a_1 _07212_ (.A1(_01705_),
    .A2(\rs2_content[26] ),
    .B1(\rs2_content[25] ),
    .B2(_01702_),
    .X(_01706_));
 sky130_fd_sc_hd__inv_2 _07213_ (.A(\rs2_content[26] ),
    .Y(_01707_));
 sky130_fd_sc_hd__o2bb2a_1 _07214_ (.A1_N(_01700_),
    .A2_N(\rs2_content[27] ),
    .B1(_01707_),
    .B2(\leorv32_alu.input1[26] ),
    .X(_01708_));
 sky130_fd_sc_hd__a21boi_1 _07215_ (.A1(_01704_),
    .A2(_01706_),
    .B1_N(_01708_),
    .Y(_01709_));
 sky130_fd_sc_hd__or2_1 _07216_ (.A(_01701_),
    .B(_01709_),
    .X(_01710_));
 sky130_fd_sc_hd__clkinv_2 _07217_ (.A(\leorv32_alu.input1[23] ),
    .Y(_01711_));
 sky130_fd_sc_hd__inv_2 _07218_ (.A(\leorv32_alu.input1[22] ),
    .Y(_01712_));
 sky130_fd_sc_hd__a22oi_1 _07219_ (.A1(_01711_),
    .A2(\rs2_content[23] ),
    .B1(\rs2_content[22] ),
    .B2(_01712_),
    .Y(_01713_));
 sky130_fd_sc_hd__clkinv_2 _07220_ (.A(\leorv32_alu.input1[21] ),
    .Y(_01714_));
 sky130_fd_sc_hd__inv_2 _07221_ (.A(\leorv32_alu.input1[20] ),
    .Y(_01715_));
 sky130_fd_sc_hd__a22oi_1 _07222_ (.A1(_01714_),
    .A2(\rs2_content[21] ),
    .B1(\rs2_content[20] ),
    .B2(_01715_),
    .Y(_01716_));
 sky130_fd_sc_hd__buf_4 _07223_ (.A(\leorv32_alu.input1[19] ),
    .X(_01717_));
 sky130_fd_sc_hd__inv_2 _07224_ (.A(\rs2_content[19] ),
    .Y(_01718_));
 sky130_fd_sc_hd__inv_2 _07225_ (.A(\rs2_content[18] ),
    .Y(_01719_));
 sky130_fd_sc_hd__o22a_1 _07226_ (.A1(\leorv32_alu.input1[19] ),
    .A2(_01718_),
    .B1(_01719_),
    .B2(\leorv32_alu.input1[18] ),
    .X(_01720_));
 sky130_fd_sc_hd__or2b_1 _07227_ (.A(\leorv32_alu.input1[17] ),
    .B_N(\rs2_content[17] ),
    .X(_01721_));
 sky130_fd_sc_hd__or2b_1 _07228_ (.A(\leorv32_alu.input1[16] ),
    .B_N(\rs2_content[16] ),
    .X(_01722_));
 sky130_fd_sc_hd__buf_4 _07229_ (.A(\leorv32_alu.input1[17] ),
    .X(_01723_));
 sky130_fd_sc_hd__and2b_1 _07230_ (.A_N(\rs2_content[17] ),
    .B(_01723_),
    .X(_01724_));
 sky130_fd_sc_hd__a221o_1 _07231_ (.A1(\leorv32_alu.input1[18] ),
    .A2(_01719_),
    .B1(_01721_),
    .B2(_01722_),
    .C1(_01724_),
    .X(_01725_));
 sky130_fd_sc_hd__nor2_1 _07232_ (.A(_01715_),
    .B(\rs2_content[20] ),
    .Y(_01726_));
 sky130_fd_sc_hd__a221o_1 _07233_ (.A1(_01717_),
    .A2(_01718_),
    .B1(_01720_),
    .B2(_01725_),
    .C1(_01726_),
    .X(_01727_));
 sky130_fd_sc_hd__nor2_1 _07234_ (.A(_01712_),
    .B(\rs2_content[22] ),
    .Y(_01728_));
 sky130_fd_sc_hd__nor2_1 _07235_ (.A(_01714_),
    .B(\rs2_content[21] ),
    .Y(_01729_));
 sky130_fd_sc_hd__a211o_1 _07236_ (.A1(_01716_),
    .A2(_01727_),
    .B1(_01728_),
    .C1(_01729_),
    .X(_01730_));
 sky130_fd_sc_hd__inv_2 _07237_ (.A(\rs2_content[24] ),
    .Y(_01731_));
 sky130_fd_sc_hd__nand2_1 _07238_ (.A(_01708_),
    .B(_01706_),
    .Y(_01732_));
 sky130_fd_sc_hd__a2111o_1 _07239_ (.A1(\leorv32_alu.input1[24] ),
    .A2(_01731_),
    .B1(_01701_),
    .C1(_01704_),
    .D1(_01732_),
    .X(_01733_));
 sky130_fd_sc_hd__nor2_1 _07240_ (.A(_01711_),
    .B(\rs2_content[23] ),
    .Y(_01734_));
 sky130_fd_sc_hd__a211o_1 _07241_ (.A1(_01713_),
    .A2(_01730_),
    .B1(_01733_),
    .C1(_01734_),
    .X(_01735_));
 sky130_fd_sc_hd__clkbuf_4 _07242_ (.A(\leorv32_alu.input1[28] ),
    .X(_01736_));
 sky130_fd_sc_hd__a21oi_1 _07243_ (.A1(_01736_),
    .A2(_01698_),
    .B1(_01697_),
    .Y(_01737_));
 sky130_fd_sc_hd__nand2_1 _07244_ (.A(_01699_),
    .B(_01737_),
    .Y(_01738_));
 sky130_fd_sc_hd__a21o_1 _07245_ (.A1(_01710_),
    .A2(_01735_),
    .B1(_01738_),
    .X(_01739_));
 sky130_fd_sc_hd__o21ai_1 _07246_ (.A1(_01697_),
    .A2(_01699_),
    .B1(_01739_),
    .Y(_01740_));
 sky130_fd_sc_hd__inv_2 _07247_ (.A(\rs2_content[15] ),
    .Y(_01741_));
 sky130_fd_sc_hd__inv_2 _07248_ (.A(\rs2_content[14] ),
    .Y(_01742_));
 sky130_fd_sc_hd__o22a_1 _07249_ (.A1(\leorv32_alu.input1[15] ),
    .A2(_01741_),
    .B1(_01742_),
    .B2(\leorv32_alu.input1[14] ),
    .X(_01743_));
 sky130_fd_sc_hd__inv_2 _07250_ (.A(\rs2_content[13] ),
    .Y(_01744_));
 sky130_fd_sc_hd__inv_2 _07251_ (.A(\rs2_content[12] ),
    .Y(_01745_));
 sky130_fd_sc_hd__o22a_1 _07252_ (.A1(\leorv32_alu.input1[13] ),
    .A2(_01744_),
    .B1(_01745_),
    .B2(\leorv32_alu.input1[12] ),
    .X(_01746_));
 sky130_fd_sc_hd__clkbuf_4 _07253_ (.A(\leorv32_alu.input1[12] ),
    .X(_01747_));
 sky130_fd_sc_hd__inv_2 _07254_ (.A(\rs2_content[11] ),
    .Y(_01748_));
 sky130_fd_sc_hd__buf_6 _07255_ (.A(\leorv32_alu.input1[11] ),
    .X(_01749_));
 sky130_fd_sc_hd__inv_2 _07256_ (.A(\rs2_content[10] ),
    .Y(_01750_));
 sky130_fd_sc_hd__inv_2 _07257_ (.A(\rs2_content[9] ),
    .Y(_01751_));
 sky130_fd_sc_hd__buf_4 _07258_ (.A(\leorv32_alu.input1[9] ),
    .X(_01752_));
 sky130_fd_sc_hd__a22o_1 _07259_ (.A1(\leorv32_alu.input1[10] ),
    .A2(_01750_),
    .B1(_01751_),
    .B2(_01752_),
    .X(_01753_));
 sky130_fd_sc_hd__clkinv_2 _07260_ (.A(\leorv32_alu.input1[8] ),
    .Y(_01754_));
 sky130_fd_sc_hd__o2bb2a_1 _07261_ (.A1_N(\rs2_content[8] ),
    .A2_N(_01754_),
    .B1(\leorv32_alu.input1[9] ),
    .B2(_01751_),
    .X(_01755_));
 sky130_fd_sc_hd__o22a_1 _07262_ (.A1(\leorv32_alu.input1[11] ),
    .A2(_01748_),
    .B1(_01750_),
    .B2(\leorv32_alu.input1[10] ),
    .X(_01756_));
 sky130_fd_sc_hd__o21a_1 _07263_ (.A1(_01753_),
    .A2(_01755_),
    .B1(_01756_),
    .X(_01757_));
 sky130_fd_sc_hd__a221o_1 _07264_ (.A1(_01747_),
    .A2(_01745_),
    .B1(_01748_),
    .B2(_01749_),
    .C1(_01757_),
    .X(_01758_));
 sky130_fd_sc_hd__a22o_1 _07265_ (.A1(\leorv32_alu.input1[14] ),
    .A2(_01742_),
    .B1(_01744_),
    .B2(\leorv32_alu.input1[13] ),
    .X(_01759_));
 sky130_fd_sc_hd__a21o_1 _07266_ (.A1(_01746_),
    .A2(_01758_),
    .B1(_01759_),
    .X(_01760_));
 sky130_fd_sc_hd__and2_1 _07267_ (.A(\leorv32_alu.input1[15] ),
    .B(_01741_),
    .X(_01761_));
 sky130_fd_sc_hd__a21o_1 _07268_ (.A1(_01743_),
    .A2(_01760_),
    .B1(_01761_),
    .X(_01762_));
 sky130_fd_sc_hd__inv_2 _07269_ (.A(\leorv32_alu.input1[5] ),
    .Y(_01763_));
 sky130_fd_sc_hd__buf_4 _07270_ (.A(\leorv32_alu.input1[4] ),
    .X(_01764_));
 sky130_fd_sc_hd__inv_2 _07271_ (.A(_01764_),
    .Y(_01765_));
 sky130_fd_sc_hd__clkinv_2 _07272_ (.A(\leorv32_alu.input1[7] ),
    .Y(_01766_));
 sky130_fd_sc_hd__inv_2 _07273_ (.A(\leorv32_alu.input1[6] ),
    .Y(_01767_));
 sky130_fd_sc_hd__a22o_1 _07274_ (.A1(_01766_),
    .A2(\rs2_content[7] ),
    .B1(\rs2_content[6] ),
    .B2(_01767_),
    .X(_01768_));
 sky130_fd_sc_hd__a221o_1 _07275_ (.A1(_01763_),
    .A2(\rs2_content[5] ),
    .B1(\rs2_content[4] ),
    .B2(_01765_),
    .C1(_01768_),
    .X(_01769_));
 sky130_fd_sc_hd__buf_6 _07276_ (.A(\rs2_content[3] ),
    .X(_01770_));
 sky130_fd_sc_hd__inv_2 _07277_ (.A(\leorv32_alu.input1[3] ),
    .Y(_01771_));
 sky130_fd_sc_hd__buf_8 _07278_ (.A(\rs2_content[2] ),
    .X(_01772_));
 sky130_fd_sc_hd__clkinv_2 _07279_ (.A(\leorv32_alu.input1[2] ),
    .Y(_01773_));
 sky130_fd_sc_hd__a22o_1 _07280_ (.A1(_01771_),
    .A2(_01770_),
    .B1(_01772_),
    .B2(_01773_),
    .X(_01774_));
 sky130_fd_sc_hd__inv_2 _07281_ (.A(\leorv32_alu.input1[1] ),
    .Y(_01775_));
 sky130_fd_sc_hd__inv_2 _07282_ (.A(\leorv32_alu.input1[0] ),
    .Y(_01776_));
 sky130_fd_sc_hd__o22a_1 _07283_ (.A1(_01775_),
    .A2(\rs2_content[1] ),
    .B1(\rs2_content[0] ),
    .B2(_01776_),
    .X(_01777_));
 sky130_fd_sc_hd__buf_4 _07284_ (.A(\leorv32_alu.input1[1] ),
    .X(_01778_));
 sky130_fd_sc_hd__clkinv_2 _07285_ (.A(\rs2_content[1] ),
    .Y(_01779_));
 sky130_fd_sc_hd__nor2_1 _07286_ (.A(_01778_),
    .B(_01779_),
    .Y(_01780_));
 sky130_fd_sc_hd__o22a_1 _07287_ (.A1(_01773_),
    .A2(_01772_),
    .B1(_01777_),
    .B2(_01780_),
    .X(_01781_));
 sky130_fd_sc_hd__or2_1 _07288_ (.A(_01774_),
    .B(_01781_),
    .X(_01782_));
 sky130_fd_sc_hd__o221a_1 _07289_ (.A1(_01765_),
    .A2(\rs2_content[4] ),
    .B1(_01770_),
    .B2(_01771_),
    .C1(_01782_),
    .X(_01783_));
 sky130_fd_sc_hd__buf_4 _07290_ (.A(\leorv32_alu.input1[7] ),
    .X(_01784_));
 sky130_fd_sc_hd__inv_2 _07291_ (.A(\rs2_content[7] ),
    .Y(_01785_));
 sky130_fd_sc_hd__inv_2 _07292_ (.A(\rs2_content[6] ),
    .Y(_01786_));
 sky130_fd_sc_hd__a2bb2o_1 _07293_ (.A1_N(\rs2_content[5] ),
    .A2_N(_01763_),
    .B1(\leorv32_alu.input1[6] ),
    .B2(_01786_),
    .X(_01787_));
 sky130_fd_sc_hd__o22a_1 _07294_ (.A1(_01784_),
    .A2(_01785_),
    .B1(_01786_),
    .B2(\leorv32_alu.input1[6] ),
    .X(_01788_));
 sky130_fd_sc_hd__or2b_1 _07295_ (.A(_01753_),
    .B_N(_01755_),
    .X(_01789_));
 sky130_fd_sc_hd__nor2_1 _07296_ (.A(_01754_),
    .B(\rs2_content[8] ),
    .Y(_01790_));
 sky130_fd_sc_hd__or3b_1 _07297_ (.A(_01761_),
    .B(_01790_),
    .C_N(_01743_),
    .X(_01791_));
 sky130_fd_sc_hd__nand2_1 _07298_ (.A(_01756_),
    .B(_01746_),
    .Y(_01792_));
 sky130_fd_sc_hd__a221o_1 _07299_ (.A1(\leorv32_alu.input1[12] ),
    .A2(_01745_),
    .B1(_01748_),
    .B2(\leorv32_alu.input1[11] ),
    .C1(_01759_),
    .X(_01793_));
 sky130_fd_sc_hd__or4_2 _07300_ (.A(_01789_),
    .B(_01791_),
    .C(_01792_),
    .D(_01793_),
    .X(_01794_));
 sky130_fd_sc_hd__a221o_1 _07301_ (.A1(_01784_),
    .A2(_01785_),
    .B1(_01787_),
    .B2(_01788_),
    .C1(_01794_),
    .X(_01795_));
 sky130_fd_sc_hd__o21bai_1 _07302_ (.A1(_01769_),
    .A2(_01783_),
    .B1_N(_01795_),
    .Y(_01796_));
 sky130_fd_sc_hd__and2_1 _07303_ (.A(_01721_),
    .B(_01722_),
    .X(_01797_));
 sky130_fd_sc_hd__nand4_1 _07304_ (.A(_01720_),
    .B(_01716_),
    .C(_01713_),
    .D(_01797_),
    .Y(_01798_));
 sky130_fd_sc_hd__inv_2 _07305_ (.A(\leorv32_alu.input1[16] ),
    .Y(_01799_));
 sky130_fd_sc_hd__a2bb2o_1 _07306_ (.A1_N(\rs2_content[16] ),
    .A2_N(_01799_),
    .B1(\leorv32_alu.input1[18] ),
    .B2(_01719_),
    .X(_01800_));
 sky130_fd_sc_hd__or4_1 _07307_ (.A(_01728_),
    .B(_01734_),
    .C(_01724_),
    .D(_01726_),
    .X(_01801_));
 sky130_fd_sc_hd__a2111o_1 _07308_ (.A1(_01717_),
    .A2(_01718_),
    .B1(_01729_),
    .C1(_01800_),
    .D1(_01801_),
    .X(_01802_));
 sky130_fd_sc_hd__or4_2 _07309_ (.A(_01738_),
    .B(_01733_),
    .C(_01798_),
    .D(_01802_),
    .X(_01803_));
 sky130_fd_sc_hd__a21oi_1 _07310_ (.A1(_01762_),
    .A2(_01796_),
    .B1(_01803_),
    .Y(_01804_));
 sky130_fd_sc_hd__nor3_1 _07311_ (.A(\leorv32_alu.input1[30] ),
    .B(_01692_),
    .C(_01695_),
    .Y(_01805_));
 sky130_fd_sc_hd__inv_2 _07312_ (.A(\rs2_content[0] ),
    .Y(_01806_));
 sky130_fd_sc_hd__clkbuf_4 _07313_ (.A(\leorv32_alu.input1[0] ),
    .X(_01807_));
 sky130_fd_sc_hd__a221o_1 _07314_ (.A1(_01778_),
    .A2(_01779_),
    .B1(_01806_),
    .B2(_01807_),
    .C1(_01774_),
    .X(_01808_));
 sky130_fd_sc_hd__a211o_1 _07315_ (.A1(_01776_),
    .A2(\rs2_content[0] ),
    .B1(_01787_),
    .C1(_01780_),
    .X(_01809_));
 sky130_fd_sc_hd__o22a_1 _07316_ (.A1(_01766_),
    .A2(\rs2_content[7] ),
    .B1(_01770_),
    .B2(_01771_),
    .X(_01810_));
 sky130_fd_sc_hd__o221a_1 _07317_ (.A1(_01765_),
    .A2(\rs2_content[4] ),
    .B1(_01772_),
    .B2(_01773_),
    .C1(_01810_),
    .X(_01811_));
 sky130_fd_sc_hd__or4b_1 _07318_ (.A(_01794_),
    .B(_01808_),
    .C(_01809_),
    .D_N(_01811_),
    .X(_01812_));
 sky130_fd_sc_hd__or3_2 _07319_ (.A(_01803_),
    .B(_01769_),
    .C(_01812_),
    .X(_01813_));
 sky130_fd_sc_hd__o41a_1 _07320_ (.A1(_01691_),
    .A2(_01740_),
    .A3(_01804_),
    .A4(_01805_),
    .B1(_01813_),
    .X(_01814_));
 sky130_fd_sc_hd__nor2_1 _07321_ (.A(_01688_),
    .B(\J_type_imm[12] ),
    .Y(_01815_));
 sky130_fd_sc_hd__nand2_4 _07322_ (.A(_01689_),
    .B(_01815_),
    .Y(_01816_));
 sky130_fd_sc_hd__nor2b_2 _07323_ (.A(\J_type_imm[13] ),
    .B_N(\J_type_imm[12] ),
    .Y(_01817_));
 sky130_fd_sc_hd__or3_1 _07324_ (.A(_01696_),
    .B(_01740_),
    .C(_01804_),
    .X(_01818_));
 sky130_fd_sc_hd__and3b_1 _07325_ (.A_N(_01691_),
    .B(_01813_),
    .C(_01818_),
    .X(_01819_));
 sky130_fd_sc_hd__and3_1 _07326_ (.A(_01687_),
    .B(_01817_),
    .C(_01819_),
    .X(_01820_));
 sky130_fd_sc_hd__o21ba_1 _07327_ (.A1(_01814_),
    .A2(_01816_),
    .B1_N(_01820_),
    .X(_01821_));
 sky130_fd_sc_hd__or2_1 _07328_ (.A(\J_type_imm[13] ),
    .B(\J_type_imm[12] ),
    .X(_01822_));
 sky130_fd_sc_hd__buf_2 _07329_ (.A(_01822_),
    .X(_01823_));
 sky130_fd_sc_hd__nor2_1 _07330_ (.A(_01687_),
    .B(_01823_),
    .Y(_01824_));
 sky130_fd_sc_hd__nand2_1 _07331_ (.A(_01813_),
    .B(_01824_),
    .Y(_01825_));
 sky130_fd_sc_hd__buf_4 _07332_ (.A(\J_type_imm[12] ),
    .X(_01826_));
 sky130_fd_sc_hd__and3_2 _07333_ (.A(_01687_),
    .B(\J_type_imm[13] ),
    .C(_01826_),
    .X(_01827_));
 sky130_fd_sc_hd__nor2_4 _07334_ (.A(\J_type_imm[13] ),
    .B(\J_type_imm[12] ),
    .Y(_01828_));
 sky130_fd_sc_hd__nand2_4 _07335_ (.A(_01687_),
    .B(_01828_),
    .Y(_01829_));
 sky130_fd_sc_hd__o2bb2a_1 _07336_ (.A1_N(_01814_),
    .A2_N(_01827_),
    .B1(_01829_),
    .B2(_01819_),
    .X(_01830_));
 sky130_fd_sc_hd__nand3_1 _07337_ (.A(_01821_),
    .B(_01825_),
    .C(_01830_),
    .Y(_01831_));
 sky130_fd_sc_hd__nand2_4 _07338_ (.A(_01688_),
    .B(_01817_),
    .Y(_01832_));
 sky130_fd_sc_hd__or2_1 _07339_ (.A(_01813_),
    .B(_01832_),
    .X(_01833_));
 sky130_fd_sc_hd__or2b_1 _07340_ (.A(_01831_),
    .B_N(_01833_),
    .X(_01834_));
 sky130_fd_sc_hd__or2_1 _07341_ (.A(_01690_),
    .B(_01834_),
    .X(_01835_));
 sky130_fd_sc_hd__buf_2 _07342_ (.A(_01835_),
    .X(_01836_));
 sky130_fd_sc_hd__clkbuf_4 _07343_ (.A(_01836_),
    .X(_01837_));
 sky130_fd_sc_hd__a21oi_1 _07344_ (.A1(_01541_),
    .A2(_01683_),
    .B1(_01837_),
    .Y(_01838_));
 sky130_fd_sc_hd__and3_1 _07345_ (.A(\PC[4] ),
    .B(\PC[3] ),
    .C(\PC[2] ),
    .X(_01839_));
 sky130_fd_sc_hd__and2_1 _07346_ (.A(\PC[5] ),
    .B(_01839_),
    .X(_01840_));
 sky130_fd_sc_hd__and3_1 _07347_ (.A(\PC[7] ),
    .B(_01591_),
    .C(_01840_),
    .X(_01841_));
 sky130_fd_sc_hd__and2_1 _07348_ (.A(\PC[8] ),
    .B(_01841_),
    .X(_01842_));
 sky130_fd_sc_hd__and3_1 _07349_ (.A(\PC[10] ),
    .B(\PC[9] ),
    .C(_01842_),
    .X(_01843_));
 sky130_fd_sc_hd__and2_1 _07350_ (.A(\PC[11] ),
    .B(_01843_),
    .X(_01844_));
 sky130_fd_sc_hd__and3_1 _07351_ (.A(\PC[13] ),
    .B(_01558_),
    .C(_01844_),
    .X(_01845_));
 sky130_fd_sc_hd__and2_1 _07352_ (.A(\PC[14] ),
    .B(_01845_),
    .X(_01846_));
 sky130_fd_sc_hd__and3_1 _07353_ (.A(\PC[16] ),
    .B(_01615_),
    .C(_01846_),
    .X(_01847_));
 sky130_fd_sc_hd__and2_1 _07354_ (.A(\PC[17] ),
    .B(_01847_),
    .X(_01848_));
 sky130_fd_sc_hd__and3_1 _07355_ (.A(\PC[19] ),
    .B(\PC[18] ),
    .C(_01848_),
    .X(_01849_));
 sky130_fd_sc_hd__and2_1 _07356_ (.A(_01546_),
    .B(_01849_),
    .X(_01850_));
 sky130_fd_sc_hd__and3_1 _07357_ (.A(\PC[22] ),
    .B(\PC[21] ),
    .C(_01850_),
    .X(_01851_));
 sky130_fd_sc_hd__xnor2_2 _07358_ (.A(\PC[23] ),
    .B(_01851_),
    .Y(_01852_));
 sky130_fd_sc_hd__and4bb_1 _07359_ (.A_N(\instr[3] ),
    .B_N(\instr[2] ),
    .C(\instr[1] ),
    .D(\instr[0] ),
    .X(_01853_));
 sky130_fd_sc_hd__clkbuf_4 _07360_ (.A(_01853_),
    .X(_01854_));
 sky130_fd_sc_hd__nand2_2 _07361_ (.A(_01531_),
    .B(_01854_),
    .Y(_01855_));
 sky130_fd_sc_hd__clkbuf_4 _07362_ (.A(_01855_),
    .X(_01856_));
 sky130_fd_sc_hd__a221oi_1 _07363_ (.A1(_01684_),
    .A2(_01838_),
    .B1(_01852_),
    .B2(_01837_),
    .C1(_01856_),
    .Y(_01857_));
 sky130_fd_sc_hd__nand4_4 _07364_ (.A(\instr[2] ),
    .B(\instr[1] ),
    .C(\instr[0] ),
    .D(_01531_),
    .Y(_01858_));
 sky130_fd_sc_hd__buf_2 _07365_ (.A(_01858_),
    .X(_01859_));
 sky130_fd_sc_hd__buf_4 _07366_ (.A(_01859_),
    .X(_01860_));
 sky130_fd_sc_hd__nor2_8 _07367_ (.A(\instr[3] ),
    .B(_01860_),
    .Y(_01861_));
 sky130_fd_sc_hd__nor2_1 _07368_ (.A(_01539_),
    .B(\leorv32_alu.input1[22] ),
    .Y(_01862_));
 sky130_fd_sc_hd__or2_1 _07369_ (.A(\leorv32_alu.input1[21] ),
    .B(\leorv32_alu.input1[20] ),
    .X(_01863_));
 sky130_fd_sc_hd__nand2_1 _07370_ (.A(_01537_),
    .B(\leorv32_alu.input1[20] ),
    .Y(_01864_));
 sky130_fd_sc_hd__or2_1 _07371_ (.A(_01537_),
    .B(\leorv32_alu.input1[20] ),
    .X(_01865_));
 sky130_fd_sc_hd__nand2_1 _07372_ (.A(_01864_),
    .B(_01865_),
    .Y(_01866_));
 sky130_fd_sc_hd__buf_4 _07373_ (.A(\leorv32_alu.input1[18] ),
    .X(_01867_));
 sky130_fd_sc_hd__clkbuf_4 _07374_ (.A(\leorv32_alu.input1[16] ),
    .X(_01868_));
 sky130_fd_sc_hd__or4_1 _07375_ (.A(_01717_),
    .B(_01867_),
    .C(_01723_),
    .D(_01868_),
    .X(_01869_));
 sky130_fd_sc_hd__buf_4 _07376_ (.A(\leorv32_alu.input1[15] ),
    .X(_01870_));
 sky130_fd_sc_hd__clkbuf_4 _07377_ (.A(\leorv32_alu.input1[14] ),
    .X(_01871_));
 sky130_fd_sc_hd__buf_4 _07378_ (.A(\leorv32_alu.input1[13] ),
    .X(_01872_));
 sky130_fd_sc_hd__or2_1 _07379_ (.A(_01872_),
    .B(_01747_),
    .X(_01873_));
 sky130_fd_sc_hd__or3_1 _07380_ (.A(_01870_),
    .B(_01871_),
    .C(_01873_),
    .X(_01874_));
 sky130_fd_sc_hd__and2_1 _07381_ (.A(_01536_),
    .B(_01874_),
    .X(_01875_));
 sky130_fd_sc_hd__xor2_4 _07382_ (.A(_01535_),
    .B(_01749_),
    .X(_01876_));
 sky130_fd_sc_hd__buf_4 _07383_ (.A(\leorv32_alu.input1[10] ),
    .X(_01877_));
 sky130_fd_sc_hd__nor2_1 _07384_ (.A(_01602_),
    .B(_01877_),
    .Y(_01878_));
 sky130_fd_sc_hd__inv_2 _07385_ (.A(\barrel_shifter_right.arith ),
    .Y(_01879_));
 sky130_fd_sc_hd__inv_2 _07386_ (.A(_01877_),
    .Y(_01880_));
 sky130_fd_sc_hd__nor2_4 _07387_ (.A(_01879_),
    .B(_01880_),
    .Y(_01881_));
 sky130_fd_sc_hd__nor2_4 _07388_ (.A(_01878_),
    .B(_01881_),
    .Y(_01882_));
 sky130_fd_sc_hd__and2_1 _07389_ (.A(_01567_),
    .B(_01752_),
    .X(_01883_));
 sky130_fd_sc_hd__or2_1 _07390_ (.A(_01567_),
    .B(_01752_),
    .X(_01884_));
 sky130_fd_sc_hd__or2b_1 _07391_ (.A(_01883_),
    .B_N(_01884_),
    .X(_01885_));
 sky130_fd_sc_hd__clkinv_2 _07392_ (.A(_01885_),
    .Y(_01886_));
 sky130_fd_sc_hd__buf_2 _07393_ (.A(\B_type_imm[7] ),
    .X(_01887_));
 sky130_fd_sc_hd__nand2_2 _07394_ (.A(_01887_),
    .B(_01784_),
    .Y(_01888_));
 sky130_fd_sc_hd__nand2_1 _07395_ (.A(_01595_),
    .B(\leorv32_alu.input1[6] ),
    .Y(_01889_));
 sky130_fd_sc_hd__clkbuf_2 _07396_ (.A(\B_type_imm[5] ),
    .X(_01890_));
 sky130_fd_sc_hd__nand2_1 _07397_ (.A(_01890_),
    .B(\leorv32_alu.input1[5] ),
    .Y(_01891_));
 sky130_fd_sc_hd__buf_2 _07398_ (.A(\I_type_imm[4] ),
    .X(_01892_));
 sky130_fd_sc_hd__nand2_1 _07399_ (.A(_01892_),
    .B(_01764_),
    .Y(_01893_));
 sky130_fd_sc_hd__inv_2 _07400_ (.A(_01893_),
    .Y(_01894_));
 sky130_fd_sc_hd__or2_1 _07401_ (.A(_01892_),
    .B(_01764_),
    .X(_01895_));
 sky130_fd_sc_hd__nand2_1 _07402_ (.A(_01893_),
    .B(_01895_),
    .Y(_01896_));
 sky130_fd_sc_hd__buf_2 _07403_ (.A(\I_type_imm[3] ),
    .X(_01897_));
 sky130_fd_sc_hd__buf_4 _07404_ (.A(\leorv32_alu.input1[3] ),
    .X(_01898_));
 sky130_fd_sc_hd__or2_1 _07405_ (.A(_01897_),
    .B(_01898_),
    .X(_01899_));
 sky130_fd_sc_hd__clkbuf_4 _07406_ (.A(\I_type_imm[2] ),
    .X(_01900_));
 sky130_fd_sc_hd__buf_4 _07407_ (.A(\leorv32_alu.input1[2] ),
    .X(_01901_));
 sky130_fd_sc_hd__nor2_1 _07408_ (.A(_01900_),
    .B(_01901_),
    .Y(_01902_));
 sky130_fd_sc_hd__nand2_2 _07409_ (.A(\I_type_imm[0] ),
    .B(\leorv32_alu.input1[0] ),
    .Y(_01903_));
 sky130_fd_sc_hd__xnor2_2 _07410_ (.A(\I_type_imm[1] ),
    .B(_01778_),
    .Y(_01904_));
 sky130_fd_sc_hd__nand2_1 _07411_ (.A(\I_type_imm[1] ),
    .B(_01778_),
    .Y(_01905_));
 sky130_fd_sc_hd__o21a_1 _07412_ (.A1(_01903_),
    .A2(_01904_),
    .B1(_01905_),
    .X(_01906_));
 sky130_fd_sc_hd__nand2_1 _07413_ (.A(_01900_),
    .B(_01901_),
    .Y(_01907_));
 sky130_fd_sc_hd__nand2_1 _07414_ (.A(_01897_),
    .B(_01898_),
    .Y(_01908_));
 sky130_fd_sc_hd__o211ai_1 _07415_ (.A1(_01902_),
    .A2(_01906_),
    .B1(_01907_),
    .C1(_01908_),
    .Y(_01909_));
 sky130_fd_sc_hd__and3b_1 _07416_ (.A_N(_01896_),
    .B(_01899_),
    .C(_01909_),
    .X(_01910_));
 sky130_fd_sc_hd__or2_1 _07417_ (.A(_01890_),
    .B(\leorv32_alu.input1[5] ),
    .X(_01911_));
 sky130_fd_sc_hd__nand2_1 _07418_ (.A(_01891_),
    .B(_01911_),
    .Y(_01912_));
 sky130_fd_sc_hd__o21bai_1 _07419_ (.A1(_01894_),
    .A2(_01910_),
    .B1_N(_01912_),
    .Y(_01913_));
 sky130_fd_sc_hd__or2_1 _07420_ (.A(_01595_),
    .B(\leorv32_alu.input1[6] ),
    .X(_01914_));
 sky130_fd_sc_hd__nand2_1 _07421_ (.A(_01889_),
    .B(_01914_),
    .Y(_01915_));
 sky130_fd_sc_hd__a21o_1 _07422_ (.A1(_01891_),
    .A2(_01913_),
    .B1(_01915_),
    .X(_01916_));
 sky130_fd_sc_hd__clkbuf_4 _07423_ (.A(\B_type_imm[8] ),
    .X(_01917_));
 sky130_fd_sc_hd__and2_1 _07424_ (.A(_01917_),
    .B(\leorv32_alu.input1[8] ),
    .X(_01918_));
 sky130_fd_sc_hd__nor2_1 _07425_ (.A(_01917_),
    .B(\leorv32_alu.input1[8] ),
    .Y(_01919_));
 sky130_fd_sc_hd__or2_2 _07426_ (.A(_01918_),
    .B(_01919_),
    .X(_01920_));
 sky130_fd_sc_hd__nor2_2 _07427_ (.A(_01887_),
    .B(_01784_),
    .Y(_01921_));
 sky130_fd_sc_hd__a311oi_4 _07428_ (.A1(_01888_),
    .A2(_01889_),
    .A3(_01916_),
    .B1(_01920_),
    .C1(_01921_),
    .Y(_01922_));
 sky130_fd_sc_hd__o221a_1 _07429_ (.A1(_01602_),
    .A2(_01877_),
    .B1(_01883_),
    .B2(_01918_),
    .C1(_01884_),
    .X(_01923_));
 sky130_fd_sc_hd__a211o_1 _07430_ (.A1(\B_type_imm[12] ),
    .A2(_01749_),
    .B1(_01923_),
    .C1(_01881_),
    .X(_01924_));
 sky130_fd_sc_hd__o21ai_1 _07431_ (.A1(_01535_),
    .A2(_01749_),
    .B1(_01924_),
    .Y(_01925_));
 sky130_fd_sc_hd__inv_2 _07432_ (.A(_01925_),
    .Y(_01926_));
 sky130_fd_sc_hd__a41oi_4 _07433_ (.A1(_01876_),
    .A2(_01882_),
    .A3(_01886_),
    .A4(_01922_),
    .B1(_01926_),
    .Y(_01927_));
 sky130_fd_sc_hd__and2_1 _07434_ (.A(\B_type_imm[12] ),
    .B(_01747_),
    .X(_01928_));
 sky130_fd_sc_hd__nor2_1 _07435_ (.A(\B_type_imm[12] ),
    .B(_01747_),
    .Y(_01929_));
 sky130_fd_sc_hd__or2_1 _07436_ (.A(_01928_),
    .B(_01929_),
    .X(_01930_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _07437_ (.A(_01930_),
    .X(_01931_));
 sky130_fd_sc_hd__xor2_4 _07438_ (.A(\B_type_imm[12] ),
    .B(_01872_),
    .X(_01932_));
 sky130_fd_sc_hd__clkinv_2 _07439_ (.A(_01932_),
    .Y(_01933_));
 sky130_fd_sc_hd__nand2_1 _07440_ (.A(_01535_),
    .B(_01871_),
    .Y(_01934_));
 sky130_fd_sc_hd__or2_1 _07441_ (.A(\B_type_imm[12] ),
    .B(_01871_),
    .X(_01935_));
 sky130_fd_sc_hd__nand2_1 _07442_ (.A(_01934_),
    .B(_01935_),
    .Y(_01936_));
 sky130_fd_sc_hd__xnor2_2 _07443_ (.A(_01535_),
    .B(_01870_),
    .Y(_01937_));
 sky130_fd_sc_hd__or4_1 _07444_ (.A(_01931_),
    .B(_01933_),
    .C(_01936_),
    .D(_01937_),
    .X(_01938_));
 sky130_fd_sc_hd__nor2_1 _07445_ (.A(_01927_),
    .B(_01938_),
    .Y(_01939_));
 sky130_fd_sc_hd__and2_1 _07446_ (.A(_01536_),
    .B(_01868_),
    .X(_01940_));
 sky130_fd_sc_hd__nor2_1 _07447_ (.A(_01536_),
    .B(_01868_),
    .Y(_01941_));
 sky130_fd_sc_hd__nor2_1 _07448_ (.A(_01940_),
    .B(_01941_),
    .Y(_01942_));
 sky130_fd_sc_hd__o21a_1 _07449_ (.A1(_01875_),
    .A2(_01939_),
    .B1(_01942_),
    .X(_01943_));
 sky130_fd_sc_hd__xor2_2 _07450_ (.A(_01536_),
    .B(_01723_),
    .X(_01944_));
 sky130_fd_sc_hd__nand2_1 _07451_ (.A(_01943_),
    .B(_01944_),
    .Y(_01945_));
 sky130_fd_sc_hd__xnor2_2 _07452_ (.A(_01536_),
    .B(_01867_),
    .Y(_01946_));
 sky130_fd_sc_hd__xor2_2 _07453_ (.A(_01536_),
    .B(_01717_),
    .X(_01947_));
 sky130_fd_sc_hd__or2b_1 _07454_ (.A(_01946_),
    .B_N(_01947_),
    .X(_01948_));
 sky130_fd_sc_hd__o2bb2a_1 _07455_ (.A1_N(_01538_),
    .A2_N(_01869_),
    .B1(_01945_),
    .B2(_01948_),
    .X(_01949_));
 sky130_fd_sc_hd__or2_1 _07456_ (.A(_01866_),
    .B(_01949_),
    .X(_01950_));
 sky130_fd_sc_hd__xnor2_2 _07457_ (.A(_01538_),
    .B(\leorv32_alu.input1[21] ),
    .Y(_01951_));
 sky130_fd_sc_hd__o2bb2a_1 _07458_ (.A1_N(_01539_),
    .A2_N(_01863_),
    .B1(_01950_),
    .B2(_01951_),
    .X(_01952_));
 sky130_fd_sc_hd__nand2_1 _07459_ (.A(_01540_),
    .B(\leorv32_alu.input1[22] ),
    .Y(_01953_));
 sky130_fd_sc_hd__o21ai_1 _07460_ (.A1(_01862_),
    .A2(_01952_),
    .B1(_01953_),
    .Y(_01954_));
 sky130_fd_sc_hd__xnor2_1 _07461_ (.A(_01540_),
    .B(\leorv32_alu.input1[23] ),
    .Y(_01955_));
 sky130_fd_sc_hd__xnor2_1 _07462_ (.A(_01954_),
    .B(_01955_),
    .Y(_01956_));
 sky130_fd_sc_hd__and2_1 _07463_ (.A(_01531_),
    .B(_01854_),
    .X(_01957_));
 sky130_fd_sc_hd__nor2_4 _07464_ (.A(_01532_),
    .B(_01957_),
    .Y(_01958_));
 sky130_fd_sc_hd__a21o_1 _07465_ (.A1(_01861_),
    .A2(_01956_),
    .B1(_01958_),
    .X(_01959_));
 sky130_fd_sc_hd__a211o_1 _07466_ (.A1(_01534_),
    .A2(_01637_),
    .B1(_01857_),
    .C1(_01959_),
    .X(_01960_));
 sky130_fd_sc_hd__a21oi_1 _07467_ (.A1(_01852_),
    .A2(_01958_),
    .B1(_01529_),
    .Y(_01961_));
 sky130_fd_sc_hd__a22o_1 _07468_ (.A1(\PC[23] ),
    .A2(_01529_),
    .B1(_01960_),
    .B2(_01961_),
    .X(_01525_));
 sky130_fd_sc_hd__and2_1 _07469_ (.A(_01539_),
    .B(\leorv32_alu.input1[22] ),
    .X(_01962_));
 sky130_fd_sc_hd__nor2_1 _07470_ (.A(_01962_),
    .B(_01862_),
    .Y(_01963_));
 sky130_fd_sc_hd__xnor2_1 _07471_ (.A(_01963_),
    .B(_01952_),
    .Y(_01964_));
 sky130_fd_sc_hd__nor2b_1 _07472_ (.A(_01635_),
    .B_N(_01542_),
    .Y(_01965_));
 sky130_fd_sc_hd__o21ai_1 _07473_ (.A1(_01634_),
    .A2(_01965_),
    .B1(_01534_),
    .Y(_01966_));
 sky130_fd_sc_hd__a21oi_1 _07474_ (.A1(_01634_),
    .A2(_01965_),
    .B1(_01966_),
    .Y(_01967_));
 sky130_fd_sc_hd__or2b_1 _07475_ (.A(_01689_),
    .B_N(_01826_),
    .X(_01968_));
 sky130_fd_sc_hd__buf_2 _07476_ (.A(_01968_),
    .X(_01969_));
 sky130_fd_sc_hd__clkbuf_4 _07477_ (.A(_01969_),
    .X(_01970_));
 sky130_fd_sc_hd__clkbuf_4 _07478_ (.A(_01816_),
    .X(_01971_));
 sky130_fd_sc_hd__clkbuf_4 _07479_ (.A(_01971_),
    .X(_01972_));
 sky130_fd_sc_hd__a21oi_1 _07480_ (.A1(\PC[21] ),
    .A2(_01850_),
    .B1(\PC[22] ),
    .Y(_01973_));
 sky130_fd_sc_hd__or2_2 _07481_ (.A(_01851_),
    .B(_01973_),
    .X(_01974_));
 sky130_fd_sc_hd__a21o_1 _07482_ (.A1(_01970_),
    .A2(_01972_),
    .B1(_01974_),
    .X(_01975_));
 sky130_fd_sc_hd__a21o_1 _07483_ (.A1(_01833_),
    .A2(_01821_),
    .B1(_01974_),
    .X(_01976_));
 sky130_fd_sc_hd__xnor2_1 _07484_ (.A(_01965_),
    .B(_01682_),
    .Y(_01977_));
 sky130_fd_sc_hd__a22o_1 _07485_ (.A1(_01837_),
    .A2(_01975_),
    .B1(_01976_),
    .B2(_01977_),
    .X(_01978_));
 sky130_fd_sc_hd__nand2_8 _07486_ (.A(_01688_),
    .B(\J_type_imm[13] ),
    .Y(_01979_));
 sky130_fd_sc_hd__a31o_1 _07487_ (.A1(_01825_),
    .A2(_01979_),
    .A3(_01830_),
    .B1(_01974_),
    .X(_01980_));
 sky130_fd_sc_hd__a21oi_1 _07488_ (.A1(_01978_),
    .A2(_01980_),
    .B1(_01856_),
    .Y(_01981_));
 sky130_fd_sc_hd__a2111o_1 _07489_ (.A1(_01861_),
    .A2(_01964_),
    .B1(_01967_),
    .C1(_01981_),
    .D1(_01958_),
    .X(_01982_));
 sky130_fd_sc_hd__a21oi_1 _07490_ (.A1(_01958_),
    .A2(_01974_),
    .B1(_01529_),
    .Y(_01983_));
 sky130_fd_sc_hd__a22o_1 _07491_ (.A1(_01529_),
    .A2(\PC[22] ),
    .B1(_01982_),
    .B2(_01983_),
    .X(_01524_));
 sky130_fd_sc_hd__clkbuf_4 _07492_ (.A(\core_state[1] ),
    .X(_01984_));
 sky130_fd_sc_hd__clkbuf_4 _07493_ (.A(_01984_),
    .X(_01985_));
 sky130_fd_sc_hd__buf_4 _07494_ (.A(_01985_),
    .X(_01986_));
 sky130_fd_sc_hd__nand2_1 _07495_ (.A(_01864_),
    .B(_01950_),
    .Y(_01987_));
 sky130_fd_sc_hd__xnor2_1 _07496_ (.A(_01951_),
    .B(_01987_),
    .Y(_01988_));
 sky130_fd_sc_hd__xnor2_1 _07497_ (.A(_01545_),
    .B(_01633_),
    .Y(_01989_));
 sky130_fd_sc_hd__nand2_1 _07498_ (.A(\instr[3] ),
    .B(_01989_),
    .Y(_01990_));
 sky130_fd_sc_hd__o211a_1 _07499_ (.A1(\instr[3] ),
    .A2(_01988_),
    .B1(_01990_),
    .C1(_01532_),
    .X(_01991_));
 sky130_fd_sc_hd__or2_1 _07500_ (.A(_01836_),
    .B(_01855_),
    .X(_01992_));
 sky130_fd_sc_hd__clkbuf_4 _07501_ (.A(_01992_),
    .X(_01993_));
 sky130_fd_sc_hd__nand2_4 _07502_ (.A(_01860_),
    .B(_01993_),
    .Y(_01994_));
 sky130_fd_sc_hd__xnor2_2 _07503_ (.A(\PC[21] ),
    .B(_01850_),
    .Y(_01995_));
 sky130_fd_sc_hd__xnor2_1 _07504_ (.A(_01545_),
    .B(_01681_),
    .Y(_01996_));
 sky130_fd_sc_hd__clkbuf_4 _07505_ (.A(_01984_),
    .X(_01997_));
 sky130_fd_sc_hd__o221ai_1 _07506_ (.A1(_01994_),
    .A2(_01995_),
    .B1(_01996_),
    .B2(_01993_),
    .C1(_01997_),
    .Y(_01998_));
 sky130_fd_sc_hd__o22a_1 _07507_ (.A1(_01986_),
    .A2(\PC[21] ),
    .B1(_01991_),
    .B2(_01998_),
    .X(_01523_));
 sky130_fd_sc_hd__xnor2_2 _07508_ (.A(_01546_),
    .B(_01849_),
    .Y(_01999_));
 sky130_fd_sc_hd__nand2_4 _07509_ (.A(\instr[3] ),
    .B(_01532_),
    .Y(_02000_));
 sky130_fd_sc_hd__and3_1 _07510_ (.A(_01548_),
    .B(_01631_),
    .C(_01638_),
    .X(_02001_));
 sky130_fd_sc_hd__a21oi_1 _07511_ (.A1(_01548_),
    .A2(_01631_),
    .B1(_01638_),
    .Y(_02002_));
 sky130_fd_sc_hd__or3_1 _07512_ (.A(_02000_),
    .B(_02001_),
    .C(_02002_),
    .X(_02003_));
 sky130_fd_sc_hd__o21ai_1 _07513_ (.A1(_01675_),
    .A2(_01679_),
    .B1(_01678_),
    .Y(_02004_));
 sky130_fd_sc_hd__and3_1 _07514_ (.A(_01638_),
    .B(_01676_),
    .C(_02004_),
    .X(_02005_));
 sky130_fd_sc_hd__a21oi_1 _07515_ (.A1(_01676_),
    .A2(_02004_),
    .B1(_01638_),
    .Y(_02006_));
 sky130_fd_sc_hd__o21a_1 _07516_ (.A1(_01972_),
    .A2(_01999_),
    .B1(_01836_),
    .X(_02007_));
 sky130_fd_sc_hd__inv_2 _07517_ (.A(_01836_),
    .Y(_02008_));
 sky130_fd_sc_hd__o32a_1 _07518_ (.A1(_02005_),
    .A2(_02006_),
    .A3(_02007_),
    .B1(_01999_),
    .B2(_02008_),
    .X(_02009_));
 sky130_fd_sc_hd__nand2_1 _07519_ (.A(_01866_),
    .B(_01949_),
    .Y(_02010_));
 sky130_fd_sc_hd__nand2_1 _07520_ (.A(_01950_),
    .B(_02010_),
    .Y(_02011_));
 sky130_fd_sc_hd__or2_1 _07521_ (.A(\instr[3] ),
    .B(_01860_),
    .X(_02012_));
 sky130_fd_sc_hd__buf_4 _07522_ (.A(_02012_),
    .X(_02013_));
 sky130_fd_sc_hd__nand2_4 _07523_ (.A(_01860_),
    .B(_01855_),
    .Y(_02014_));
 sky130_fd_sc_hd__o221a_1 _07524_ (.A1(_01856_),
    .A2(_02009_),
    .B1(_02011_),
    .B2(_02013_),
    .C1(_02014_),
    .X(_02015_));
 sky130_fd_sc_hd__a221o_1 _07525_ (.A1(_01958_),
    .A2(_01999_),
    .B1(_02003_),
    .B2(_02015_),
    .C1(_01529_),
    .X(_02016_));
 sky130_fd_sc_hd__a21bo_1 _07526_ (.A1(_01529_),
    .A2(_01546_),
    .B1_N(_02016_),
    .X(_01522_));
 sky130_fd_sc_hd__a21oi_1 _07527_ (.A1(\PC[18] ),
    .A2(_01848_),
    .B1(\PC[19] ),
    .Y(_02017_));
 sky130_fd_sc_hd__or2_1 _07528_ (.A(_01849_),
    .B(_02017_),
    .X(_02018_));
 sky130_fd_sc_hd__o21ai_1 _07529_ (.A1(_01994_),
    .A2(_02018_),
    .B1(_01997_),
    .Y(_02019_));
 sky130_fd_sc_hd__a211o_1 _07530_ (.A1(_01548_),
    .A2(_01629_),
    .B1(_01549_),
    .C1(_01628_),
    .X(_02020_));
 sky130_fd_sc_hd__nor2_2 _07531_ (.A(_01837_),
    .B(_01855_),
    .Y(_02021_));
 sky130_fd_sc_hd__or3_1 _07532_ (.A(_01675_),
    .B(_01678_),
    .C(_01679_),
    .X(_02022_));
 sky130_fd_sc_hd__o21ai_1 _07533_ (.A1(_01723_),
    .A2(_01868_),
    .B1(_01539_),
    .Y(_02023_));
 sky130_fd_sc_hd__a21oi_1 _07534_ (.A1(_01945_),
    .A2(_02023_),
    .B1(_01946_),
    .Y(_02024_));
 sky130_fd_sc_hd__a21oi_1 _07535_ (.A1(_01540_),
    .A2(_01867_),
    .B1(_02024_),
    .Y(_02025_));
 sky130_fd_sc_hd__xnor2_1 _07536_ (.A(_01947_),
    .B(_02025_),
    .Y(_02026_));
 sky130_fd_sc_hd__a32o_1 _07537_ (.A1(_02021_),
    .A2(_02004_),
    .A3(_02022_),
    .B1(_02026_),
    .B2(_01861_),
    .X(_02027_));
 sky130_fd_sc_hd__a31o_1 _07538_ (.A1(_01631_),
    .A2(_01534_),
    .A3(_02020_),
    .B1(_02027_),
    .X(_02028_));
 sky130_fd_sc_hd__o22a_1 _07539_ (.A1(_01997_),
    .A2(\PC[19] ),
    .B1(_02019_),
    .B2(_02028_),
    .X(_01521_));
 sky130_fd_sc_hd__xnor2_2 _07540_ (.A(\PC[18] ),
    .B(_01848_),
    .Y(_02029_));
 sky130_fd_sc_hd__o21a_1 _07541_ (.A1(_02014_),
    .A2(_02029_),
    .B1(_01997_),
    .X(_02030_));
 sky130_fd_sc_hd__nand3_1 _07542_ (.A(_01945_),
    .B(_01946_),
    .C(_02023_),
    .Y(_02031_));
 sky130_fd_sc_hd__and2b_1 _07543_ (.A_N(_02024_),
    .B(_02031_),
    .X(_02032_));
 sky130_fd_sc_hd__o21ai_1 _07544_ (.A1(_01551_),
    .A2(_01627_),
    .B1(_01534_),
    .Y(_02033_));
 sky130_fd_sc_hd__nor2_1 _07545_ (.A(_01628_),
    .B(_02033_),
    .Y(_02034_));
 sky130_fd_sc_hd__and2_1 _07546_ (.A(_01979_),
    .B(_02029_),
    .X(_02035_));
 sky130_fd_sc_hd__nand2_1 _07547_ (.A(\PC[17] ),
    .B(_01540_),
    .Y(_02036_));
 sky130_fd_sc_hd__a21oi_1 _07548_ (.A1(_02036_),
    .A2(_01674_),
    .B1(_01640_),
    .Y(_02037_));
 sky130_fd_sc_hd__a31o_1 _07549_ (.A1(_01640_),
    .A2(_02036_),
    .A3(_01674_),
    .B1(_01836_),
    .X(_02038_));
 sky130_fd_sc_hd__o22a_1 _07550_ (.A1(_02008_),
    .A2(_02035_),
    .B1(_02037_),
    .B2(_02038_),
    .X(_02039_));
 sky130_fd_sc_hd__a211oi_1 _07551_ (.A1(_01690_),
    .A2(_02029_),
    .B1(_02039_),
    .C1(_01856_),
    .Y(_02040_));
 sky130_fd_sc_hd__a211oi_1 _07552_ (.A1(_01861_),
    .A2(_02032_),
    .B1(_02034_),
    .C1(_02040_),
    .Y(_02041_));
 sky130_fd_sc_hd__o2bb2a_1 _07553_ (.A1_N(_02030_),
    .A2_N(_02041_),
    .B1(_01986_),
    .B2(\PC[18] ),
    .X(_01520_));
 sky130_fd_sc_hd__nor2_1 _07554_ (.A(\PC[17] ),
    .B(_01847_),
    .Y(_02042_));
 sky130_fd_sc_hd__or2_1 _07555_ (.A(_01848_),
    .B(_02042_),
    .X(_02043_));
 sky130_fd_sc_hd__o2111a_1 _07556_ (.A1(_01673_),
    .A2(_01672_),
    .B1(_01669_),
    .C1(_01670_),
    .D1(_01671_),
    .X(_02044_));
 sky130_fd_sc_hd__or3b_1 _07557_ (.A(_01837_),
    .B(_02044_),
    .C_N(_01674_),
    .X(_02045_));
 sky130_fd_sc_hd__o21a_1 _07558_ (.A1(_02008_),
    .A2(_02043_),
    .B1(_02045_),
    .X(_02046_));
 sky130_fd_sc_hd__nor2_1 _07559_ (.A(_01856_),
    .B(_02046_),
    .Y(_02047_));
 sky130_fd_sc_hd__or2_1 _07560_ (.A(_01940_),
    .B(_01943_),
    .X(_02048_));
 sky130_fd_sc_hd__xnor2_1 _07561_ (.A(_01944_),
    .B(_02048_),
    .Y(_02049_));
 sky130_fd_sc_hd__nor2_1 _07562_ (.A(_02013_),
    .B(_02049_),
    .Y(_02050_));
 sky130_fd_sc_hd__nand2_1 _07563_ (.A(_01554_),
    .B(_01625_),
    .Y(_02051_));
 sky130_fd_sc_hd__o21ai_1 _07564_ (.A1(_02014_),
    .A2(_02043_),
    .B1(_01984_),
    .Y(_02052_));
 sky130_fd_sc_hd__a31o_1 _07565_ (.A1(_01626_),
    .A2(_01534_),
    .A3(_02051_),
    .B1(_02052_),
    .X(_02053_));
 sky130_fd_sc_hd__o32a_1 _07566_ (.A1(_02047_),
    .A2(_02050_),
    .A3(_02053_),
    .B1(\PC[17] ),
    .B2(_01986_),
    .X(_01519_));
 sky130_fd_sc_hd__nand2_1 _07567_ (.A(_01615_),
    .B(_01846_),
    .Y(_02054_));
 sky130_fd_sc_hd__xor2_2 _07568_ (.A(\PC[16] ),
    .B(_02054_),
    .X(_02055_));
 sky130_fd_sc_hd__o21a_1 _07569_ (.A1(_01832_),
    .A2(_02055_),
    .B1(_01837_),
    .X(_02056_));
 sky130_fd_sc_hd__a21oi_1 _07570_ (.A1(_01666_),
    .A2(_01670_),
    .B1(_01668_),
    .Y(_02057_));
 sky130_fd_sc_hd__a21oi_1 _07571_ (.A1(_01615_),
    .A2(_01540_),
    .B1(_02057_),
    .Y(_02058_));
 sky130_fd_sc_hd__xnor2_1 _07572_ (.A(_01667_),
    .B(_02058_),
    .Y(_02059_));
 sky130_fd_sc_hd__o22a_1 _07573_ (.A1(_02008_),
    .A2(_02055_),
    .B1(_02056_),
    .B2(_02059_),
    .X(_02060_));
 sky130_fd_sc_hd__nor2_1 _07574_ (.A(_01856_),
    .B(_02060_),
    .Y(_02061_));
 sky130_fd_sc_hd__or3_1 _07575_ (.A(_01942_),
    .B(_01875_),
    .C(_01939_),
    .X(_02062_));
 sky130_fd_sc_hd__or2b_1 _07576_ (.A(_01943_),
    .B_N(_02062_),
    .X(_02063_));
 sky130_fd_sc_hd__o221ai_1 _07577_ (.A1(_02014_),
    .A2(_02055_),
    .B1(_02063_),
    .B2(_02013_),
    .C1(_01997_),
    .Y(_02064_));
 sky130_fd_sc_hd__a21o_1 _07578_ (.A1(_01611_),
    .A2(_01622_),
    .B1(_01613_),
    .X(_02065_));
 sky130_fd_sc_hd__or2_1 _07579_ (.A(_01618_),
    .B(_02065_),
    .X(_02066_));
 sky130_fd_sc_hd__nand2_1 _07580_ (.A(_01616_),
    .B(_02066_),
    .Y(_02067_));
 sky130_fd_sc_hd__a21oi_1 _07581_ (.A1(_01557_),
    .A2(_02067_),
    .B1(_02000_),
    .Y(_02068_));
 sky130_fd_sc_hd__o21a_1 _07582_ (.A1(_01557_),
    .A2(_02067_),
    .B1(_02068_),
    .X(_02069_));
 sky130_fd_sc_hd__o32a_1 _07583_ (.A1(_02061_),
    .A2(_02064_),
    .A3(_02069_),
    .B1(\PC[16] ),
    .B2(_01986_),
    .X(_01518_));
 sky130_fd_sc_hd__or2_1 _07584_ (.A(_01615_),
    .B(_01846_),
    .X(_02070_));
 sky130_fd_sc_hd__nand2_2 _07585_ (.A(_02054_),
    .B(_02070_),
    .Y(_02071_));
 sky130_fd_sc_hd__o21a_1 _07586_ (.A1(_01972_),
    .A2(_02071_),
    .B1(_01837_),
    .X(_02072_));
 sky130_fd_sc_hd__and3_1 _07587_ (.A(_01666_),
    .B(_01668_),
    .C(_01670_),
    .X(_02073_));
 sky130_fd_sc_hd__or2_1 _07588_ (.A(_02057_),
    .B(_02073_),
    .X(_02074_));
 sky130_fd_sc_hd__o221a_1 _07589_ (.A1(_01833_),
    .A2(_02071_),
    .B1(_02072_),
    .B2(_02074_),
    .C1(_01979_),
    .X(_02075_));
 sky130_fd_sc_hd__a211o_1 _07590_ (.A1(_01690_),
    .A2(_02071_),
    .B1(_02075_),
    .C1(_01856_),
    .X(_02076_));
 sky130_fd_sc_hd__nor2_1 _07591_ (.A(_01927_),
    .B(_01931_),
    .Y(_02077_));
 sky130_fd_sc_hd__a22o_1 _07592_ (.A1(_01540_),
    .A2(_01873_),
    .B1(_01932_),
    .B2(_02077_),
    .X(_02078_));
 sky130_fd_sc_hd__a21boi_1 _07593_ (.A1(_01935_),
    .A2(_02078_),
    .B1_N(_01934_),
    .Y(_02079_));
 sky130_fd_sc_hd__xnor2_1 _07594_ (.A(_01937_),
    .B(_02079_),
    .Y(_02080_));
 sky130_fd_sc_hd__nand2_1 _07595_ (.A(_01618_),
    .B(_02065_),
    .Y(_02081_));
 sky130_fd_sc_hd__nand2_1 _07596_ (.A(_02066_),
    .B(_02081_),
    .Y(_02082_));
 sky130_fd_sc_hd__xnor2_2 _07597_ (.A(_01558_),
    .B(_01844_),
    .Y(_02083_));
 sky130_fd_sc_hd__a21oi_1 _07598_ (.A1(_01690_),
    .A2(_02083_),
    .B1(_01855_),
    .Y(_02084_));
 sky130_fd_sc_hd__a21oi_1 _07599_ (.A1(_01831_),
    .A2(_02084_),
    .B1(_01958_),
    .Y(_02085_));
 sky130_fd_sc_hd__o221a_1 _07600_ (.A1(_02000_),
    .A2(_02082_),
    .B1(_02085_),
    .B2(_02071_),
    .C1(_01984_),
    .X(_02086_));
 sky130_fd_sc_hd__o21a_1 _07601_ (.A1(_02013_),
    .A2(_02080_),
    .B1(_02086_),
    .X(_02087_));
 sky130_fd_sc_hd__o2bb2a_1 _07602_ (.A1_N(_02076_),
    .A2_N(_02087_),
    .B1(_01986_),
    .B2(_01615_),
    .X(_01517_));
 sky130_fd_sc_hd__nor2_1 _07603_ (.A(\PC[14] ),
    .B(_01845_),
    .Y(_02088_));
 sky130_fd_sc_hd__or2_2 _07604_ (.A(_01846_),
    .B(_02088_),
    .X(_02089_));
 sky130_fd_sc_hd__a21o_1 _07605_ (.A1(_01958_),
    .A2(_02089_),
    .B1(_01529_),
    .X(_02090_));
 sky130_fd_sc_hd__a21o_1 _07606_ (.A1(_01979_),
    .A2(_02089_),
    .B1(_02008_),
    .X(_02091_));
 sky130_fd_sc_hd__a21o_1 _07607_ (.A1(_01832_),
    .A2(_01972_),
    .B1(_02089_),
    .X(_02092_));
 sky130_fd_sc_hd__and3_1 _07608_ (.A(_01641_),
    .B(_01662_),
    .C(_01665_),
    .X(_02093_));
 sky130_fd_sc_hd__a21oi_1 _07609_ (.A1(_01662_),
    .A2(_01665_),
    .B1(_01641_),
    .Y(_02094_));
 sky130_fd_sc_hd__a211o_1 _07610_ (.A1(_01837_),
    .A2(_02092_),
    .B1(_02093_),
    .C1(_02094_),
    .X(_02095_));
 sky130_fd_sc_hd__a22o_1 _07611_ (.A1(_01690_),
    .A2(_02089_),
    .B1(_02091_),
    .B2(_02095_),
    .X(_02096_));
 sky130_fd_sc_hd__xor2_1 _07612_ (.A(_01936_),
    .B(_02078_),
    .X(_02097_));
 sky130_fd_sc_hd__nor2_1 _07613_ (.A(_01621_),
    .B(_01561_),
    .Y(_02098_));
 sky130_fd_sc_hd__a21oi_1 _07614_ (.A1(_01611_),
    .A2(_02098_),
    .B1(_01614_),
    .Y(_02099_));
 sky130_fd_sc_hd__a31o_1 _07615_ (.A1(_01611_),
    .A2(_01614_),
    .A3(_02098_),
    .B1(_02000_),
    .X(_02100_));
 sky130_fd_sc_hd__o22a_1 _07616_ (.A1(_02013_),
    .A2(_02097_),
    .B1(_02099_),
    .B2(_02100_),
    .X(_02101_));
 sky130_fd_sc_hd__o211a_1 _07617_ (.A1(_01856_),
    .A2(_02096_),
    .B1(_02101_),
    .C1(_02014_),
    .X(_02102_));
 sky130_fd_sc_hd__a2bb2o_1 _07618_ (.A1_N(_02090_),
    .A2_N(_02102_),
    .B1(\PC[14] ),
    .B2(_01529_),
    .X(_01516_));
 sky130_fd_sc_hd__nor2_1 _07619_ (.A(_01928_),
    .B(_02077_),
    .Y(_02103_));
 sky130_fd_sc_hd__xnor2_1 _07620_ (.A(_01932_),
    .B(_02103_),
    .Y(_02104_));
 sky130_fd_sc_hd__and2_1 _07621_ (.A(_01861_),
    .B(_02104_),
    .X(_02105_));
 sky130_fd_sc_hd__nor2_1 _07622_ (.A(_01563_),
    .B(_01610_),
    .Y(_02106_));
 sky130_fd_sc_hd__or2_1 _07623_ (.A(_01559_),
    .B(_01560_),
    .X(_02107_));
 sky130_fd_sc_hd__o211a_1 _07624_ (.A1(_02106_),
    .A2(_02107_),
    .B1(_01611_),
    .C1(_01562_),
    .X(_02108_));
 sky130_fd_sc_hd__a21oi_1 _07625_ (.A1(_01558_),
    .A2(_01844_),
    .B1(\PC[13] ),
    .Y(_02109_));
 sky130_fd_sc_hd__or2_1 _07626_ (.A(_01845_),
    .B(_02109_),
    .X(_02110_));
 sky130_fd_sc_hd__nor2_1 _07627_ (.A(_01994_),
    .B(_02110_),
    .Y(_02111_));
 sky130_fd_sc_hd__a211o_1 _07628_ (.A1(_01534_),
    .A2(_02108_),
    .B1(_02111_),
    .C1(_01528_),
    .X(_02112_));
 sky130_fd_sc_hd__or2_1 _07629_ (.A(_01661_),
    .B(_01664_),
    .X(_02113_));
 sky130_fd_sc_hd__and3_1 _07630_ (.A(_01665_),
    .B(_02021_),
    .C(_02113_),
    .X(_02114_));
 sky130_fd_sc_hd__o32a_1 _07631_ (.A1(_02105_),
    .A2(_02112_),
    .A3(_02114_),
    .B1(\PC[13] ),
    .B2(_01986_),
    .X(_01515_));
 sky130_fd_sc_hd__or2_1 _07632_ (.A(_01559_),
    .B(_01563_),
    .X(_02115_));
 sky130_fd_sc_hd__xnor2_1 _07633_ (.A(_01610_),
    .B(_02115_),
    .Y(_02116_));
 sky130_fd_sc_hd__a21o_1 _07634_ (.A1(_01643_),
    .A2(_01657_),
    .B1(_01659_),
    .X(_02117_));
 sky130_fd_sc_hd__xor2_1 _07635_ (.A(_01558_),
    .B(_01539_),
    .X(_02118_));
 sky130_fd_sc_hd__xnor2_1 _07636_ (.A(_02117_),
    .B(_02118_),
    .Y(_02119_));
 sky130_fd_sc_hd__o221ai_1 _07637_ (.A1(_01833_),
    .A2(_02083_),
    .B1(_02119_),
    .B2(_01836_),
    .C1(_01979_),
    .Y(_02120_));
 sky130_fd_sc_hd__nand2_1 _07638_ (.A(_01927_),
    .B(_01931_),
    .Y(_02121_));
 sky130_fd_sc_hd__or2b_1 _07639_ (.A(_02077_),
    .B_N(_02121_),
    .X(_02122_));
 sky130_fd_sc_hd__o2bb2a_1 _07640_ (.A1_N(_02084_),
    .A2_N(_02120_),
    .B1(_02122_),
    .B2(_02012_),
    .X(_02123_));
 sky130_fd_sc_hd__o221ai_1 _07641_ (.A1(_02083_),
    .A2(_02085_),
    .B1(_02116_),
    .B2(_02000_),
    .C1(_02123_),
    .Y(_02124_));
 sky130_fd_sc_hd__mux2_1 _07642_ (.A0(_01558_),
    .A1(_02124_),
    .S(_01985_),
    .X(_02125_));
 sky130_fd_sc_hd__clkbuf_1 _07643_ (.A(_02125_),
    .X(_01514_));
 sky130_fd_sc_hd__nand2_1 _07644_ (.A(_01658_),
    .B(_01643_),
    .Y(_02126_));
 sky130_fd_sc_hd__xor2_1 _07645_ (.A(_02126_),
    .B(_01657_),
    .X(_02127_));
 sky130_fd_sc_hd__nor2_1 _07646_ (.A(\PC[11] ),
    .B(_01843_),
    .Y(_02128_));
 sky130_fd_sc_hd__or2_1 _07647_ (.A(_01844_),
    .B(_02128_),
    .X(_02129_));
 sky130_fd_sc_hd__mux2_1 _07648_ (.A0(_02127_),
    .A1(_02129_),
    .S(_01837_),
    .X(_02130_));
 sky130_fd_sc_hd__nor2_1 _07649_ (.A(_01856_),
    .B(_02130_),
    .Y(_02131_));
 sky130_fd_sc_hd__o31a_1 _07650_ (.A1(_01883_),
    .A2(_01918_),
    .A3(_01922_),
    .B1(_01884_),
    .X(_02132_));
 sky130_fd_sc_hd__a21oi_1 _07651_ (.A1(_01882_),
    .A2(_02132_),
    .B1(_01881_),
    .Y(_02133_));
 sky130_fd_sc_hd__xor2_1 _07652_ (.A(_01876_),
    .B(_02133_),
    .X(_02134_));
 sky130_fd_sc_hd__o21a_1 _07653_ (.A1(_01565_),
    .A2(_01609_),
    .B1(_01608_),
    .X(_02135_));
 sky130_fd_sc_hd__o31ai_1 _07654_ (.A1(_01565_),
    .A2(_01609_),
    .A3(_01608_),
    .B1(_01534_),
    .Y(_02136_));
 sky130_fd_sc_hd__o221a_1 _07655_ (.A1(_02014_),
    .A2(_02129_),
    .B1(_02135_),
    .B2(_02136_),
    .C1(_01985_),
    .X(_02137_));
 sky130_fd_sc_hd__o21ai_1 _07656_ (.A1(_02013_),
    .A2(_02134_),
    .B1(_02137_),
    .Y(_02138_));
 sky130_fd_sc_hd__o22a_1 _07657_ (.A1(_01997_),
    .A2(\PC[11] ),
    .B1(_02131_),
    .B2(_02138_),
    .X(_01513_));
 sky130_fd_sc_hd__a21oi_1 _07658_ (.A1(\PC[9] ),
    .A2(_01842_),
    .B1(\PC[10] ),
    .Y(_02139_));
 sky130_fd_sc_hd__nor2_2 _07659_ (.A(_01843_),
    .B(_02139_),
    .Y(_02140_));
 sky130_fd_sc_hd__o21ba_1 _07660_ (.A1(_01570_),
    .A2(_01656_),
    .B1_N(_01566_),
    .X(_02141_));
 sky130_fd_sc_hd__xnor2_1 _07661_ (.A(_01605_),
    .B(_02141_),
    .Y(_02142_));
 sky130_fd_sc_hd__nor2_1 _07662_ (.A(_01836_),
    .B(_02142_),
    .Y(_02143_));
 sky130_fd_sc_hd__a211o_1 _07663_ (.A1(_01834_),
    .A2(_02140_),
    .B1(_02143_),
    .C1(_01690_),
    .X(_02144_));
 sky130_fd_sc_hd__o21a_1 _07664_ (.A1(_01979_),
    .A2(_02140_),
    .B1(_01957_),
    .X(_02145_));
 sky130_fd_sc_hd__xor2_1 _07665_ (.A(_01882_),
    .B(_02132_),
    .X(_02146_));
 sky130_fd_sc_hd__o21ba_1 _07666_ (.A1(_01570_),
    .A2(_01600_),
    .B1_N(_01566_),
    .X(_02147_));
 sky130_fd_sc_hd__xnor2_1 _07667_ (.A(_02147_),
    .B(_01604_),
    .Y(_02148_));
 sky130_fd_sc_hd__a22o_1 _07668_ (.A1(_01861_),
    .A2(_02146_),
    .B1(_02148_),
    .B2(_01533_),
    .X(_02149_));
 sky130_fd_sc_hd__a221o_1 _07669_ (.A1(_01958_),
    .A2(_02140_),
    .B1(_02144_),
    .B2(_02145_),
    .C1(_02149_),
    .X(_02150_));
 sky130_fd_sc_hd__mux2_1 _07670_ (.A0(\PC[10] ),
    .A1(_02150_),
    .S(_01985_),
    .X(_02151_));
 sky130_fd_sc_hd__clkbuf_1 _07671_ (.A(_02151_),
    .X(_01512_));
 sky130_fd_sc_hd__xnor2_2 _07672_ (.A(\PC[9] ),
    .B(_01842_),
    .Y(_02152_));
 sky130_fd_sc_hd__o21ai_1 _07673_ (.A1(_02014_),
    .A2(_02152_),
    .B1(_01997_),
    .Y(_02153_));
 sky130_fd_sc_hd__nor2_1 _07674_ (.A(_01918_),
    .B(_01922_),
    .Y(_02154_));
 sky130_fd_sc_hd__xnor2_1 _07675_ (.A(_01886_),
    .B(_02154_),
    .Y(_02155_));
 sky130_fd_sc_hd__xor2_1 _07676_ (.A(_01570_),
    .B(_01600_),
    .X(_02156_));
 sky130_fd_sc_hd__xnor2_1 _07677_ (.A(_01570_),
    .B(_01656_),
    .Y(_02157_));
 sky130_fd_sc_hd__mux2_1 _07678_ (.A0(_02157_),
    .A1(_02152_),
    .S(_01837_),
    .X(_02158_));
 sky130_fd_sc_hd__nor2_1 _07679_ (.A(_01856_),
    .B(_02158_),
    .Y(_02159_));
 sky130_fd_sc_hd__a221o_1 _07680_ (.A1(_01861_),
    .A2(_02155_),
    .B1(_02156_),
    .B2(_01534_),
    .C1(_02159_),
    .X(_02160_));
 sky130_fd_sc_hd__o22a_1 _07681_ (.A1(_01997_),
    .A2(\PC[9] ),
    .B1(_02153_),
    .B2(_02160_),
    .X(_01511_));
 sky130_fd_sc_hd__nor2_1 _07682_ (.A(\PC[8] ),
    .B(_01841_),
    .Y(_02161_));
 sky130_fd_sc_hd__nor2_2 _07683_ (.A(_01842_),
    .B(_02161_),
    .Y(_02162_));
 sky130_fd_sc_hd__or2_1 _07684_ (.A(_01644_),
    .B(_01654_),
    .X(_02163_));
 sky130_fd_sc_hd__a21oi_1 _07685_ (.A1(_01597_),
    .A2(_02163_),
    .B1(_01577_),
    .Y(_02164_));
 sky130_fd_sc_hd__nor2_1 _07686_ (.A(_01575_),
    .B(_02164_),
    .Y(_02165_));
 sky130_fd_sc_hd__xnor2_1 _07687_ (.A(_01573_),
    .B(_02165_),
    .Y(_02166_));
 sky130_fd_sc_hd__nor2_1 _07688_ (.A(_01836_),
    .B(_02166_),
    .Y(_02167_));
 sky130_fd_sc_hd__a211o_1 _07689_ (.A1(_01834_),
    .A2(_02162_),
    .B1(_02167_),
    .C1(_01690_),
    .X(_02168_));
 sky130_fd_sc_hd__o211a_1 _07690_ (.A1(_01979_),
    .A2(_02162_),
    .B1(_02168_),
    .C1(_01957_),
    .X(_02169_));
 sky130_fd_sc_hd__and2_1 _07691_ (.A(_01571_),
    .B(_01572_),
    .X(_02170_));
 sky130_fd_sc_hd__nand2_1 _07692_ (.A(_01589_),
    .B(_01594_),
    .Y(_02171_));
 sky130_fd_sc_hd__a21oi_1 _07693_ (.A1(_01597_),
    .A2(_02171_),
    .B1(_01577_),
    .Y(_02172_));
 sky130_fd_sc_hd__or3_1 _07694_ (.A(_01575_),
    .B(_02170_),
    .C(_02172_),
    .X(_02173_));
 sky130_fd_sc_hd__o21ai_1 _07695_ (.A1(_01575_),
    .A2(_02172_),
    .B1(_02170_),
    .Y(_02174_));
 sky130_fd_sc_hd__and2_1 _07696_ (.A(_01889_),
    .B(_01916_),
    .X(_02175_));
 sky130_fd_sc_hd__o211a_1 _07697_ (.A1(_01921_),
    .A2(_02175_),
    .B1(_01920_),
    .C1(_01888_),
    .X(_02176_));
 sky130_fd_sc_hd__nor2_1 _07698_ (.A(_01922_),
    .B(_02176_),
    .Y(_02177_));
 sky130_fd_sc_hd__a32o_1 _07699_ (.A1(_01533_),
    .A2(_02173_),
    .A3(_02174_),
    .B1(_01861_),
    .B2(_02177_),
    .X(_02178_));
 sky130_fd_sc_hd__a211o_1 _07700_ (.A1(_01958_),
    .A2(_02162_),
    .B1(_02169_),
    .C1(_02178_),
    .X(_02179_));
 sky130_fd_sc_hd__mux2_1 _07701_ (.A0(\PC[8] ),
    .A1(_02179_),
    .S(_01985_),
    .X(_02180_));
 sky130_fd_sc_hd__clkbuf_1 _07702_ (.A(_02180_),
    .X(_01510_));
 sky130_fd_sc_hd__a31o_1 _07703_ (.A1(_01597_),
    .A2(_01577_),
    .A3(_02163_),
    .B1(_01993_),
    .X(_02181_));
 sky130_fd_sc_hd__a21oi_1 _07704_ (.A1(_01591_),
    .A2(_01840_),
    .B1(\PC[7] ),
    .Y(_02182_));
 sky130_fd_sc_hd__or2_1 _07705_ (.A(_01841_),
    .B(_02182_),
    .X(_02183_));
 sky130_fd_sc_hd__inv_2 _07706_ (.A(_01888_),
    .Y(_02184_));
 sky130_fd_sc_hd__nor2_1 _07707_ (.A(_02184_),
    .B(_01921_),
    .Y(_02185_));
 sky130_fd_sc_hd__xor2_1 _07708_ (.A(_02175_),
    .B(_02185_),
    .X(_02186_));
 sky130_fd_sc_hd__and3_1 _07709_ (.A(_01597_),
    .B(_01577_),
    .C(_02171_),
    .X(_02187_));
 sky130_fd_sc_hd__or3_1 _07710_ (.A(_02000_),
    .B(_02172_),
    .C(_02187_),
    .X(_02188_));
 sky130_fd_sc_hd__o221a_1 _07711_ (.A1(_01994_),
    .A2(_02183_),
    .B1(_02186_),
    .B2(_02013_),
    .C1(_02188_),
    .X(_02189_));
 sky130_fd_sc_hd__o211a_1 _07712_ (.A1(_02164_),
    .A2(_02181_),
    .B1(_02189_),
    .C1(_01985_),
    .X(_02190_));
 sky130_fd_sc_hd__o21ba_1 _07713_ (.A1(_01986_),
    .A2(\PC[7] ),
    .B1_N(_02190_),
    .X(_01509_));
 sky130_fd_sc_hd__xnor2_1 _07714_ (.A(_01591_),
    .B(_01840_),
    .Y(_02191_));
 sky130_fd_sc_hd__nor2_1 _07715_ (.A(_01994_),
    .B(_02191_),
    .Y(_02192_));
 sky130_fd_sc_hd__a21bo_1 _07716_ (.A1(_01590_),
    .A2(_01654_),
    .B1_N(_01593_),
    .X(_02193_));
 sky130_fd_sc_hd__xor2_1 _07717_ (.A(_01592_),
    .B(_02193_),
    .X(_02194_));
 sky130_fd_sc_hd__nand3_1 _07718_ (.A(_01915_),
    .B(_01891_),
    .C(_01913_),
    .Y(_02195_));
 sky130_fd_sc_hd__nand2_1 _07719_ (.A(_01916_),
    .B(_02195_),
    .Y(_02196_));
 sky130_fd_sc_hd__nand2_1 _07720_ (.A(_01590_),
    .B(_01593_),
    .Y(_02197_));
 sky130_fd_sc_hd__and2_1 _07721_ (.A(_01581_),
    .B(_01587_),
    .X(_02198_));
 sky130_fd_sc_hd__a21oi_2 _07722_ (.A1(_01579_),
    .A2(_02198_),
    .B1(_01588_),
    .Y(_02199_));
 sky130_fd_sc_hd__o21ai_1 _07723_ (.A1(_02197_),
    .A2(_02199_),
    .B1(_01590_),
    .Y(_02200_));
 sky130_fd_sc_hd__xnor2_1 _07724_ (.A(_01592_),
    .B(_02200_),
    .Y(_02201_));
 sky130_fd_sc_hd__o221a_1 _07725_ (.A1(_02013_),
    .A2(_02196_),
    .B1(_02201_),
    .B2(_02000_),
    .C1(_01985_),
    .X(_02202_));
 sky130_fd_sc_hd__o21ai_1 _07726_ (.A1(_01993_),
    .A2(_02194_),
    .B1(_02202_),
    .Y(_02203_));
 sky130_fd_sc_hd__o22a_1 _07727_ (.A1(_01997_),
    .A2(_01591_),
    .B1(_02192_),
    .B2(_02203_),
    .X(_01508_));
 sky130_fd_sc_hd__xnor2_1 _07728_ (.A(_02197_),
    .B(_01654_),
    .Y(_02204_));
 sky130_fd_sc_hd__nor2_1 _07729_ (.A(\PC[5] ),
    .B(_01839_),
    .Y(_02205_));
 sky130_fd_sc_hd__or2_1 _07730_ (.A(_01840_),
    .B(_02205_),
    .X(_02206_));
 sky130_fd_sc_hd__a211o_1 _07731_ (.A1(_01891_),
    .A2(_01911_),
    .B1(_01894_),
    .C1(_01910_),
    .X(_02207_));
 sky130_fd_sc_hd__nand2_1 _07732_ (.A(_01913_),
    .B(_02207_),
    .Y(_02208_));
 sky130_fd_sc_hd__nor2_1 _07733_ (.A(_02197_),
    .B(_02199_),
    .Y(_02209_));
 sky130_fd_sc_hd__and2_1 _07734_ (.A(_02197_),
    .B(_02199_),
    .X(_02210_));
 sky130_fd_sc_hd__or3_1 _07735_ (.A(_02209_),
    .B(_02000_),
    .C(_02210_),
    .X(_02211_));
 sky130_fd_sc_hd__o221a_1 _07736_ (.A1(_01994_),
    .A2(_02206_),
    .B1(_02208_),
    .B2(_02013_),
    .C1(_02211_),
    .X(_02212_));
 sky130_fd_sc_hd__o211a_1 _07737_ (.A1(_01993_),
    .A2(_02204_),
    .B1(_02212_),
    .C1(_01985_),
    .X(_02213_));
 sky130_fd_sc_hd__o21ba_1 _07738_ (.A1(_01986_),
    .A2(\PC[5] ),
    .B1_N(_02213_),
    .X(_01507_));
 sky130_fd_sc_hd__a21oi_1 _07739_ (.A1(\PC[3] ),
    .A2(_01585_),
    .B1(\PC[4] ),
    .Y(_02214_));
 sky130_fd_sc_hd__or2_1 _07740_ (.A(_01839_),
    .B(_02214_),
    .X(_02215_));
 sky130_fd_sc_hd__nor2_1 _07741_ (.A(_01994_),
    .B(_02215_),
    .Y(_02216_));
 sky130_fd_sc_hd__or2b_1 _07742_ (.A(_01645_),
    .B_N(_01653_),
    .X(_02217_));
 sky130_fd_sc_hd__nor3_1 _07743_ (.A(_01646_),
    .B(_01652_),
    .C(_02217_),
    .Y(_02218_));
 sky130_fd_sc_hd__o21a_1 _07744_ (.A1(_01646_),
    .A2(_01652_),
    .B1(_02217_),
    .X(_02219_));
 sky130_fd_sc_hd__and2_1 _07745_ (.A(_01899_),
    .B(_01909_),
    .X(_02220_));
 sky130_fd_sc_hd__xor2_1 _07746_ (.A(_01896_),
    .B(_02220_),
    .X(_02221_));
 sky130_fd_sc_hd__nor2_1 _07747_ (.A(\PC[4] ),
    .B(_01892_),
    .Y(_02222_));
 sky130_fd_sc_hd__nor2_1 _07748_ (.A(_02222_),
    .B(_01588_),
    .Y(_02223_));
 sky130_fd_sc_hd__xnor2_1 _07749_ (.A(_02198_),
    .B(_02223_),
    .Y(_02224_));
 sky130_fd_sc_hd__o221a_1 _07750_ (.A1(_02013_),
    .A2(_02221_),
    .B1(_02224_),
    .B2(_02000_),
    .C1(_01985_),
    .X(_02225_));
 sky130_fd_sc_hd__o31ai_1 _07751_ (.A1(_01993_),
    .A2(_02218_),
    .A3(_02219_),
    .B1(_02225_),
    .Y(_02226_));
 sky130_fd_sc_hd__o22a_1 _07752_ (.A1(_01997_),
    .A2(\PC[4] ),
    .B1(_02216_),
    .B2(_02226_),
    .X(_01506_));
 sky130_fd_sc_hd__xnor2_1 _07753_ (.A(\PC[3] ),
    .B(_01585_),
    .Y(_02227_));
 sky130_fd_sc_hd__nor2_1 _07754_ (.A(_01994_),
    .B(_02227_),
    .Y(_02228_));
 sky130_fd_sc_hd__o21a_1 _07755_ (.A1(_01647_),
    .A2(_01649_),
    .B1(_01651_),
    .X(_02229_));
 sky130_fd_sc_hd__or2b_1 _07756_ (.A(_01646_),
    .B_N(_01650_),
    .X(_02230_));
 sky130_fd_sc_hd__xnor2_1 _07757_ (.A(_02229_),
    .B(_02230_),
    .Y(_02231_));
 sky130_fd_sc_hd__nor2_1 _07758_ (.A(_01993_),
    .B(_02231_),
    .Y(_02232_));
 sky130_fd_sc_hd__o21ai_1 _07759_ (.A1(_01902_),
    .A2(_01906_),
    .B1(_01907_),
    .Y(_02233_));
 sky130_fd_sc_hd__nand2_1 _07760_ (.A(_01899_),
    .B(_01908_),
    .Y(_02234_));
 sky130_fd_sc_hd__xnor2_1 _07761_ (.A(_02233_),
    .B(_02234_),
    .Y(_02235_));
 sky130_fd_sc_hd__a21oi_1 _07762_ (.A1(_01582_),
    .A2(_01583_),
    .B1(_01586_),
    .Y(_02236_));
 sky130_fd_sc_hd__or3_1 _07763_ (.A(_01580_),
    .B(_01584_),
    .C(_02236_),
    .X(_02237_));
 sky130_fd_sc_hd__o21ai_1 _07764_ (.A1(_01580_),
    .A2(_01584_),
    .B1(_02236_),
    .Y(_02238_));
 sky130_fd_sc_hd__and3_1 _07765_ (.A(_01534_),
    .B(_02237_),
    .C(_02238_),
    .X(_02239_));
 sky130_fd_sc_hd__a211o_1 _07766_ (.A1(_01861_),
    .A2(_02235_),
    .B1(_02239_),
    .C1(_01529_),
    .X(_02240_));
 sky130_fd_sc_hd__o32a_1 _07767_ (.A1(_02228_),
    .A2(_02232_),
    .A3(_02240_),
    .B1(\PC[3] ),
    .B2(_01986_),
    .X(_01505_));
 sky130_fd_sc_hd__buf_4 _07768_ (.A(\B_type_imm[2] ),
    .X(_02241_));
 sky130_fd_sc_hd__or2_1 _07769_ (.A(_01585_),
    .B(_02241_),
    .X(_02242_));
 sky130_fd_sc_hd__and3b_1 _07770_ (.A_N(_01649_),
    .B(_02242_),
    .C(_01651_),
    .X(_02243_));
 sky130_fd_sc_hd__a21boi_1 _07771_ (.A1(_01651_),
    .A2(_02242_),
    .B1_N(_01649_),
    .Y(_02244_));
 sky130_fd_sc_hd__and2b_1 _07772_ (.A_N(_01902_),
    .B(_01907_),
    .X(_02245_));
 sky130_fd_sc_hd__xor2_1 _07773_ (.A(_01906_),
    .B(_02245_),
    .X(_02246_));
 sky130_fd_sc_hd__xnor2_1 _07774_ (.A(_01582_),
    .B(_01583_),
    .Y(_02247_));
 sky130_fd_sc_hd__o221a_1 _07775_ (.A1(_02012_),
    .A2(_02246_),
    .B1(_02247_),
    .B2(_02000_),
    .C1(_01984_),
    .X(_02248_));
 sky130_fd_sc_hd__o31a_1 _07776_ (.A1(_02243_),
    .A2(_01993_),
    .A3(_02244_),
    .B1(_02248_),
    .X(_02249_));
 sky130_fd_sc_hd__o21ai_1 _07777_ (.A1(_01585_),
    .A2(_01994_),
    .B1(_02249_),
    .Y(_02250_));
 sky130_fd_sc_hd__o21a_1 _07778_ (.A1(_01986_),
    .A2(_01585_),
    .B1(_02250_),
    .X(_01504_));
 sky130_fd_sc_hd__or2b_2 _07779_ (.A(net1),
    .B_N(\core_state[2] ),
    .X(_02251_));
 sky130_fd_sc_hd__inv_6 _07780_ (.A(_02251_),
    .Y(_02252_));
 sky130_fd_sc_hd__buf_6 _07781_ (.A(_02252_),
    .X(_02253_));
 sky130_fd_sc_hd__buf_4 _07782_ (.A(_02253_),
    .X(_02254_));
 sky130_fd_sc_hd__buf_4 _07783_ (.A(_02254_),
    .X(_00001_));
 sky130_fd_sc_hd__buf_4 _07784_ (.A(_02252_),
    .X(_02255_));
 sky130_fd_sc_hd__mux2_1 _07785_ (.A0(_01540_),
    .A1(net26),
    .S(_02255_),
    .X(_02256_));
 sky130_fd_sc_hd__clkbuf_1 _07786_ (.A(_02256_),
    .X(_01471_));
 sky130_fd_sc_hd__mux2_1 _07787_ (.A0(_01602_),
    .A1(net25),
    .S(_02255_),
    .X(_02257_));
 sky130_fd_sc_hd__clkbuf_1 _07788_ (.A(_02257_),
    .X(_01470_));
 sky130_fd_sc_hd__mux2_1 _07789_ (.A0(_01567_),
    .A1(net23),
    .S(_02255_),
    .X(_02258_));
 sky130_fd_sc_hd__clkbuf_1 _07790_ (.A(_02258_),
    .X(_01469_));
 sky130_fd_sc_hd__mux2_1 _07791_ (.A0(_01917_),
    .A1(net22),
    .S(_02255_),
    .X(_02259_));
 sky130_fd_sc_hd__clkbuf_1 _07792_ (.A(_02259_),
    .X(_01468_));
 sky130_fd_sc_hd__mux2_1 _07793_ (.A0(_01887_),
    .A1(net21),
    .S(_02255_),
    .X(_02260_));
 sky130_fd_sc_hd__clkbuf_1 _07794_ (.A(_02260_),
    .X(_01467_));
 sky130_fd_sc_hd__mux2_1 _07795_ (.A0(_01595_),
    .A1(net20),
    .S(_02255_),
    .X(_02261_));
 sky130_fd_sc_hd__clkbuf_1 _07796_ (.A(_02261_),
    .X(_01466_));
 sky130_fd_sc_hd__mux2_1 _07797_ (.A0(_01890_),
    .A1(net19),
    .S(_02255_),
    .X(_02262_));
 sky130_fd_sc_hd__clkbuf_1 _07798_ (.A(_02262_),
    .X(_01465_));
 sky130_fd_sc_hd__clkinv_4 _07799_ (.A(net18),
    .Y(_02263_));
 sky130_fd_sc_hd__buf_8 _07800_ (.A(_02263_),
    .X(_02264_));
 sky130_fd_sc_hd__nand2_8 _07801_ (.A(_02264_),
    .B(_02252_),
    .Y(_02265_));
 sky130_fd_sc_hd__buf_4 _07802_ (.A(_02265_),
    .X(_02266_));
 sky130_fd_sc_hd__o21a_1 _07803_ (.A1(_01892_),
    .A2(_00001_),
    .B1(_02266_),
    .X(_01464_));
 sky130_fd_sc_hd__buf_6 _07804_ (.A(net17),
    .X(_02267_));
 sky130_fd_sc_hd__buf_6 _07805_ (.A(_02267_),
    .X(_02268_));
 sky130_fd_sc_hd__clkbuf_4 _07806_ (.A(_02253_),
    .X(_02269_));
 sky130_fd_sc_hd__mux2_1 _07807_ (.A0(_01897_),
    .A1(_02268_),
    .S(_02269_),
    .X(_02270_));
 sky130_fd_sc_hd__clkbuf_1 _07808_ (.A(_02270_),
    .X(_01463_));
 sky130_fd_sc_hd__buf_6 _07809_ (.A(net16),
    .X(_02271_));
 sky130_fd_sc_hd__buf_8 _07810_ (.A(_02271_),
    .X(_02272_));
 sky130_fd_sc_hd__buf_8 _07811_ (.A(_02272_),
    .X(_02273_));
 sky130_fd_sc_hd__mux2_1 _07812_ (.A0(_01900_),
    .A1(_02273_),
    .S(_02269_),
    .X(_02274_));
 sky130_fd_sc_hd__clkbuf_1 _07813_ (.A(_02274_),
    .X(_01462_));
 sky130_fd_sc_hd__buf_2 _07814_ (.A(\I_type_imm[1] ),
    .X(_02275_));
 sky130_fd_sc_hd__buf_8 _07815_ (.A(net15),
    .X(_02276_));
 sky130_fd_sc_hd__buf_6 _07816_ (.A(_02276_),
    .X(_02277_));
 sky130_fd_sc_hd__clkbuf_8 _07817_ (.A(_02277_),
    .X(_02278_));
 sky130_fd_sc_hd__mux2_1 _07818_ (.A0(_02275_),
    .A1(_02278_),
    .S(_02269_),
    .X(_02279_));
 sky130_fd_sc_hd__clkbuf_1 _07819_ (.A(_02279_),
    .X(_01461_));
 sky130_fd_sc_hd__buf_8 _07820_ (.A(net14),
    .X(_02280_));
 sky130_fd_sc_hd__buf_8 _07821_ (.A(_02280_),
    .X(_02281_));
 sky130_fd_sc_hd__clkbuf_16 _07822_ (.A(_02281_),
    .X(_02282_));
 sky130_fd_sc_hd__buf_8 _07823_ (.A(_02282_),
    .X(_02283_));
 sky130_fd_sc_hd__mux2_1 _07824_ (.A0(_01564_),
    .A1(_02283_),
    .S(_02269_),
    .X(_02284_));
 sky130_fd_sc_hd__clkbuf_1 _07825_ (.A(_02284_),
    .X(_01460_));
 sky130_fd_sc_hd__inv_2 _07826_ (.A(net12),
    .Y(_02285_));
 sky130_fd_sc_hd__buf_6 _07827_ (.A(_02285_),
    .X(_02286_));
 sky130_fd_sc_hd__nand2_1 _07828_ (.A(_02286_),
    .B(_02253_),
    .Y(_02287_));
 sky130_fd_sc_hd__clkbuf_4 _07829_ (.A(_02287_),
    .X(_02288_));
 sky130_fd_sc_hd__o21a_1 _07830_ (.A1(\J_type_imm[19] ),
    .A2(_00001_),
    .B1(_02288_),
    .X(_01459_));
 sky130_fd_sc_hd__buf_4 _07831_ (.A(net11),
    .X(_02289_));
 sky130_fd_sc_hd__clkbuf_8 _07832_ (.A(_02289_),
    .X(_02290_));
 sky130_fd_sc_hd__buf_4 _07833_ (.A(_02290_),
    .X(_02291_));
 sky130_fd_sc_hd__mux2_1 _07834_ (.A0(\J_type_imm[18] ),
    .A1(_02291_),
    .S(_02269_),
    .X(_02292_));
 sky130_fd_sc_hd__clkbuf_1 _07835_ (.A(_02292_),
    .X(_01458_));
 sky130_fd_sc_hd__buf_4 _07836_ (.A(net10),
    .X(_02293_));
 sky130_fd_sc_hd__buf_6 _07837_ (.A(_02293_),
    .X(_02294_));
 sky130_fd_sc_hd__buf_6 _07838_ (.A(_02294_),
    .X(_02295_));
 sky130_fd_sc_hd__mux2_1 _07839_ (.A0(\J_type_imm[17] ),
    .A1(_02295_),
    .S(_02269_),
    .X(_02296_));
 sky130_fd_sc_hd__clkbuf_1 _07840_ (.A(_02296_),
    .X(_01457_));
 sky130_fd_sc_hd__buf_6 _07841_ (.A(net9),
    .X(_02297_));
 sky130_fd_sc_hd__buf_8 _07842_ (.A(_02297_),
    .X(_02298_));
 sky130_fd_sc_hd__buf_4 _07843_ (.A(_02298_),
    .X(_02299_));
 sky130_fd_sc_hd__mux2_1 _07844_ (.A0(\J_type_imm[16] ),
    .A1(_02299_),
    .S(_02269_),
    .X(_02300_));
 sky130_fd_sc_hd__clkbuf_1 _07845_ (.A(_02300_),
    .X(_01456_));
 sky130_fd_sc_hd__buf_4 _07846_ (.A(net8),
    .X(_02301_));
 sky130_fd_sc_hd__clkbuf_8 _07847_ (.A(_02301_),
    .X(_02302_));
 sky130_fd_sc_hd__buf_8 _07848_ (.A(_02302_),
    .X(_02303_));
 sky130_fd_sc_hd__buf_6 _07849_ (.A(_02303_),
    .X(_02304_));
 sky130_fd_sc_hd__mux2_1 _07850_ (.A0(\J_type_imm[15] ),
    .A1(_02304_),
    .S(_02269_),
    .X(_02305_));
 sky130_fd_sc_hd__clkbuf_1 _07851_ (.A(_02305_),
    .X(_01455_));
 sky130_fd_sc_hd__clkbuf_4 _07852_ (.A(_01687_),
    .X(_02306_));
 sky130_fd_sc_hd__clkbuf_4 _07853_ (.A(_02306_),
    .X(_02307_));
 sky130_fd_sc_hd__buf_4 _07854_ (.A(_02307_),
    .X(_02308_));
 sky130_fd_sc_hd__mux2_1 _07855_ (.A0(_02308_),
    .A1(net7),
    .S(_02269_),
    .X(_02309_));
 sky130_fd_sc_hd__clkbuf_1 _07856_ (.A(_02309_),
    .X(_01454_));
 sky130_fd_sc_hd__mux2_1 _07857_ (.A0(_01689_),
    .A1(net6),
    .S(_02269_),
    .X(_02310_));
 sky130_fd_sc_hd__clkbuf_1 _07858_ (.A(_02310_),
    .X(_01453_));
 sky130_fd_sc_hd__clkbuf_4 _07859_ (.A(_02252_),
    .X(_02311_));
 sky130_fd_sc_hd__mux2_1 _07860_ (.A0(_01826_),
    .A1(net5),
    .S(_02311_),
    .X(_02312_));
 sky130_fd_sc_hd__clkbuf_1 _07861_ (.A(_02312_),
    .X(_01452_));
 sky130_fd_sc_hd__buf_4 _07862_ (.A(\B_type_imm[4] ),
    .X(_02313_));
 sky130_fd_sc_hd__mux2_1 _07863_ (.A0(_02313_),
    .A1(net4),
    .S(_02311_),
    .X(_02314_));
 sky130_fd_sc_hd__clkbuf_1 _07864_ (.A(_02314_),
    .X(_01451_));
 sky130_fd_sc_hd__buf_4 _07865_ (.A(\B_type_imm[3] ),
    .X(_02315_));
 sky130_fd_sc_hd__mux2_1 _07866_ (.A0(_02315_),
    .A1(net3),
    .S(_02311_),
    .X(_02316_));
 sky130_fd_sc_hd__clkbuf_1 _07867_ (.A(_02316_),
    .X(_01450_));
 sky130_fd_sc_hd__mux2_1 _07868_ (.A0(_02241_),
    .A1(net33),
    .S(_02311_),
    .X(_02317_));
 sky130_fd_sc_hd__clkbuf_1 _07869_ (.A(_02317_),
    .X(_01449_));
 sky130_fd_sc_hd__mux2_1 _07870_ (.A0(_01648_),
    .A1(net32),
    .S(_02311_),
    .X(_02318_));
 sky130_fd_sc_hd__clkbuf_1 _07871_ (.A(_02318_),
    .X(_01448_));
 sky130_fd_sc_hd__mux2_1 _07872_ (.A0(_01642_),
    .A1(net31),
    .S(_02311_),
    .X(_02319_));
 sky130_fd_sc_hd__clkbuf_1 _07873_ (.A(_02319_),
    .X(_01447_));
 sky130_fd_sc_hd__mux2_1 _07874_ (.A0(\instr[6] ),
    .A1(net30),
    .S(_02311_),
    .X(_02320_));
 sky130_fd_sc_hd__clkbuf_1 _07875_ (.A(_02320_),
    .X(_01446_));
 sky130_fd_sc_hd__mux2_1 _07876_ (.A0(\instr[5] ),
    .A1(net29),
    .S(_02311_),
    .X(_02321_));
 sky130_fd_sc_hd__clkbuf_1 _07877_ (.A(_02321_),
    .X(_01445_));
 sky130_fd_sc_hd__mux2_1 _07878_ (.A0(_01530_),
    .A1(net28),
    .S(_02311_),
    .X(_02322_));
 sky130_fd_sc_hd__clkbuf_1 _07879_ (.A(_02322_),
    .X(_01444_));
 sky130_fd_sc_hd__mux2_1 _07880_ (.A0(\instr[3] ),
    .A1(net27),
    .S(_02311_),
    .X(_02323_));
 sky130_fd_sc_hd__clkbuf_1 _07881_ (.A(_02323_),
    .X(_01443_));
 sky130_fd_sc_hd__buf_4 _07882_ (.A(_02252_),
    .X(_02324_));
 sky130_fd_sc_hd__mux2_1 _07883_ (.A0(\instr[2] ),
    .A1(net24),
    .S(_02324_),
    .X(_02325_));
 sky130_fd_sc_hd__clkbuf_1 _07884_ (.A(_02325_),
    .X(_01442_));
 sky130_fd_sc_hd__mux2_1 _07885_ (.A0(\instr[1] ),
    .A1(net13),
    .S(_02324_),
    .X(_02326_));
 sky130_fd_sc_hd__clkbuf_1 _07886_ (.A(_02326_),
    .X(_01441_));
 sky130_fd_sc_hd__mux2_1 _07887_ (.A0(\instr[0] ),
    .A1(net2),
    .S(_02324_),
    .X(_02327_));
 sky130_fd_sc_hd__clkbuf_1 _07888_ (.A(_02327_),
    .X(_01440_));
 sky130_fd_sc_hd__clkbuf_4 _07889_ (.A(_02255_),
    .X(_02328_));
 sky130_fd_sc_hd__inv_2 _07890_ (.A(net10),
    .Y(_02329_));
 sky130_fd_sc_hd__buf_6 _07891_ (.A(_02329_),
    .X(_02330_));
 sky130_fd_sc_hd__buf_6 _07892_ (.A(_02330_),
    .X(_02331_));
 sky130_fd_sc_hd__buf_8 _07893_ (.A(net8),
    .X(_02332_));
 sky130_fd_sc_hd__buf_6 _07894_ (.A(_02332_),
    .X(_02333_));
 sky130_fd_sc_hd__buf_6 _07895_ (.A(_02333_),
    .X(_02334_));
 sky130_fd_sc_hd__buf_6 _07896_ (.A(net9),
    .X(_02335_));
 sky130_fd_sc_hd__buf_6 _07897_ (.A(_02335_),
    .X(_02336_));
 sky130_fd_sc_hd__buf_6 _07898_ (.A(_02336_),
    .X(_02337_));
 sky130_fd_sc_hd__mux4_1 _07899_ (.A0(\regs[12][31] ),
    .A1(\regs[13][31] ),
    .A2(\regs[14][31] ),
    .A3(\regs[15][31] ),
    .S0(_02334_),
    .S1(_02337_),
    .X(_02338_));
 sky130_fd_sc_hd__or2_1 _07900_ (.A(_02331_),
    .B(_02338_),
    .X(_02339_));
 sky130_fd_sc_hd__buf_8 _07901_ (.A(_02332_),
    .X(_02340_));
 sky130_fd_sc_hd__buf_12 _07902_ (.A(_02340_),
    .X(_02341_));
 sky130_fd_sc_hd__buf_6 _07903_ (.A(net9),
    .X(_02342_));
 sky130_fd_sc_hd__buf_8 _07904_ (.A(_02342_),
    .X(_02343_));
 sky130_fd_sc_hd__buf_8 _07905_ (.A(_02343_),
    .X(_02344_));
 sky130_fd_sc_hd__mux4_1 _07906_ (.A0(\regs[8][31] ),
    .A1(\regs[9][31] ),
    .A2(\regs[10][31] ),
    .A3(\regs[11][31] ),
    .S0(_02341_),
    .S1(_02344_),
    .X(_02345_));
 sky130_fd_sc_hd__clkbuf_8 _07907_ (.A(_02289_),
    .X(_02346_));
 sky130_fd_sc_hd__o21a_1 _07908_ (.A1(_02295_),
    .A2(_02345_),
    .B1(_02346_),
    .X(_02347_));
 sky130_fd_sc_hd__buf_8 _07909_ (.A(net8),
    .X(_02348_));
 sky130_fd_sc_hd__buf_6 _07910_ (.A(_02348_),
    .X(_02349_));
 sky130_fd_sc_hd__buf_8 _07911_ (.A(_02349_),
    .X(_02350_));
 sky130_fd_sc_hd__buf_6 _07912_ (.A(_02335_),
    .X(_02351_));
 sky130_fd_sc_hd__buf_6 _07913_ (.A(_02351_),
    .X(_02352_));
 sky130_fd_sc_hd__mux4_1 _07914_ (.A0(\regs[0][31] ),
    .A1(\regs[1][31] ),
    .A2(\regs[2][31] ),
    .A3(\regs[3][31] ),
    .S0(_02350_),
    .S1(_02352_),
    .X(_02353_));
 sky130_fd_sc_hd__buf_8 _07915_ (.A(_02301_),
    .X(_02354_));
 sky130_fd_sc_hd__buf_8 _07916_ (.A(_02354_),
    .X(_02355_));
 sky130_fd_sc_hd__buf_6 _07917_ (.A(_02351_),
    .X(_02356_));
 sky130_fd_sc_hd__mux4_1 _07918_ (.A0(\regs[4][31] ),
    .A1(\regs[5][31] ),
    .A2(\regs[6][31] ),
    .A3(\regs[7][31] ),
    .S0(_02355_),
    .S1(_02356_),
    .X(_02357_));
 sky130_fd_sc_hd__buf_6 _07919_ (.A(net10),
    .X(_02358_));
 sky130_fd_sc_hd__buf_8 _07920_ (.A(_02358_),
    .X(_02359_));
 sky130_fd_sc_hd__mux2_1 _07921_ (.A0(_02353_),
    .A1(_02357_),
    .S(_02359_),
    .X(_02360_));
 sky130_fd_sc_hd__inv_6 _07922_ (.A(net11),
    .Y(_02361_));
 sky130_fd_sc_hd__buf_6 _07923_ (.A(_02361_),
    .X(_02362_));
 sky130_fd_sc_hd__buf_4 _07924_ (.A(_02362_),
    .X(_02363_));
 sky130_fd_sc_hd__a22o_1 _07925_ (.A1(_02339_),
    .A2(_02347_),
    .B1(_02360_),
    .B2(_02363_),
    .X(_02364_));
 sky130_fd_sc_hd__buf_6 _07926_ (.A(_02361_),
    .X(_02365_));
 sky130_fd_sc_hd__buf_4 _07927_ (.A(_02365_),
    .X(_02366_));
 sky130_fd_sc_hd__clkbuf_8 _07928_ (.A(net9),
    .X(_02367_));
 sky130_fd_sc_hd__buf_6 _07929_ (.A(_02367_),
    .X(_02368_));
 sky130_fd_sc_hd__buf_6 _07930_ (.A(_02368_),
    .X(_02369_));
 sky130_fd_sc_hd__mux4_1 _07931_ (.A0(\regs[16][31] ),
    .A1(\regs[17][31] ),
    .A2(\regs[18][31] ),
    .A3(\regs[19][31] ),
    .S0(_02304_),
    .S1(_02369_),
    .X(_02370_));
 sky130_fd_sc_hd__buf_8 _07932_ (.A(_02302_),
    .X(_02371_));
 sky130_fd_sc_hd__buf_6 _07933_ (.A(_02371_),
    .X(_02372_));
 sky130_fd_sc_hd__clkbuf_8 _07934_ (.A(_02368_),
    .X(_02373_));
 sky130_fd_sc_hd__mux4_1 _07935_ (.A0(\regs[20][31] ),
    .A1(\regs[21][31] ),
    .A2(\regs[22][31] ),
    .A3(\regs[23][31] ),
    .S0(_02372_),
    .S1(_02373_),
    .X(_02374_));
 sky130_fd_sc_hd__buf_6 _07936_ (.A(_02293_),
    .X(_02375_));
 sky130_fd_sc_hd__buf_6 _07937_ (.A(_02375_),
    .X(_02376_));
 sky130_fd_sc_hd__mux2_1 _07938_ (.A0(_02370_),
    .A1(_02374_),
    .S(_02376_),
    .X(_02377_));
 sky130_fd_sc_hd__buf_6 _07939_ (.A(_02340_),
    .X(_02378_));
 sky130_fd_sc_hd__or2b_1 _07940_ (.A(\regs[27][31] ),
    .B_N(_02378_),
    .X(_02379_));
 sky130_fd_sc_hd__clkbuf_4 _07941_ (.A(_02301_),
    .X(_02380_));
 sky130_fd_sc_hd__clkbuf_4 _07942_ (.A(_02380_),
    .X(_02381_));
 sky130_fd_sc_hd__buf_6 _07943_ (.A(_02297_),
    .X(_02382_));
 sky130_fd_sc_hd__o21a_1 _07944_ (.A1(_02381_),
    .A2(\regs[26][31] ),
    .B1(_02382_),
    .X(_02383_));
 sky130_fd_sc_hd__buf_4 _07945_ (.A(_02354_),
    .X(_02384_));
 sky130_fd_sc_hd__mux2_1 _07946_ (.A0(\regs[24][31] ),
    .A1(\regs[25][31] ),
    .S(_02384_),
    .X(_02385_));
 sky130_fd_sc_hd__inv_2 _07947_ (.A(net9),
    .Y(_02386_));
 sky130_fd_sc_hd__buf_4 _07948_ (.A(_02386_),
    .X(_02387_));
 sky130_fd_sc_hd__buf_4 _07949_ (.A(_02387_),
    .X(_02388_));
 sky130_fd_sc_hd__buf_4 _07950_ (.A(_02388_),
    .X(_02389_));
 sky130_fd_sc_hd__buf_12 _07951_ (.A(_02358_),
    .X(_02390_));
 sky130_fd_sc_hd__a221o_1 _07952_ (.A1(_02379_),
    .A2(_02383_),
    .B1(_02385_),
    .B2(_02389_),
    .C1(_02390_),
    .X(_02391_));
 sky130_fd_sc_hd__buf_8 _07953_ (.A(_02349_),
    .X(_02392_));
 sky130_fd_sc_hd__mux2_1 _07954_ (.A0(\regs[30][31] ),
    .A1(\regs[31][31] ),
    .S(_02392_),
    .X(_02393_));
 sky130_fd_sc_hd__clkbuf_8 _07955_ (.A(_02387_),
    .X(_02394_));
 sky130_fd_sc_hd__buf_6 _07956_ (.A(_02348_),
    .X(_02395_));
 sky130_fd_sc_hd__mux2_1 _07957_ (.A0(\regs[28][31] ),
    .A1(\regs[29][31] ),
    .S(_02395_),
    .X(_02396_));
 sky130_fd_sc_hd__a21o_1 _07958_ (.A1(_02394_),
    .A2(_02396_),
    .B1(_02330_),
    .X(_02397_));
 sky130_fd_sc_hd__a21o_1 _07959_ (.A1(_02299_),
    .A2(_02393_),
    .B1(_02397_),
    .X(_02398_));
 sky130_fd_sc_hd__nand2_4 _07960_ (.A(net12),
    .B(_02252_),
    .Y(_02399_));
 sky130_fd_sc_hd__a31o_1 _07961_ (.A1(_02291_),
    .A2(_02391_),
    .A3(_02398_),
    .B1(_02399_),
    .X(_02400_));
 sky130_fd_sc_hd__a21o_1 _07962_ (.A1(_02366_),
    .A2(_02377_),
    .B1(_02400_),
    .X(_02401_));
 sky130_fd_sc_hd__o221a_1 _07963_ (.A1(\leorv32_alu.input1[31] ),
    .A2(_02328_),
    .B1(_02288_),
    .B2(_02364_),
    .C1(_02401_),
    .X(_01439_));
 sky130_fd_sc_hd__buf_6 _07964_ (.A(net9),
    .X(_02402_));
 sky130_fd_sc_hd__buf_4 _07965_ (.A(_02301_),
    .X(_02403_));
 sky130_fd_sc_hd__mux2_1 _07966_ (.A0(\regs[30][30] ),
    .A1(\regs[31][30] ),
    .S(_02403_),
    .X(_02404_));
 sky130_fd_sc_hd__and2_1 _07967_ (.A(_02402_),
    .B(_02404_),
    .X(_02405_));
 sky130_fd_sc_hd__buf_6 _07968_ (.A(_02301_),
    .X(_02406_));
 sky130_fd_sc_hd__mux2_1 _07969_ (.A0(\regs[28][30] ),
    .A1(\regs[29][30] ),
    .S(_02406_),
    .X(_02407_));
 sky130_fd_sc_hd__buf_4 _07970_ (.A(_02329_),
    .X(_02408_));
 sky130_fd_sc_hd__a21o_1 _07971_ (.A1(_02388_),
    .A2(_02407_),
    .B1(_02408_),
    .X(_02409_));
 sky130_fd_sc_hd__or2b_1 _07972_ (.A(\regs[27][30] ),
    .B_N(_02380_),
    .X(_02410_));
 sky130_fd_sc_hd__o21a_1 _07973_ (.A1(_02380_),
    .A2(\regs[26][30] ),
    .B1(_02342_),
    .X(_02411_));
 sky130_fd_sc_hd__mux2_1 _07974_ (.A0(\regs[24][30] ),
    .A1(\regs[25][30] ),
    .S(_02302_),
    .X(_02412_));
 sky130_fd_sc_hd__buf_4 _07975_ (.A(_02387_),
    .X(_02413_));
 sky130_fd_sc_hd__buf_6 _07976_ (.A(net10),
    .X(_02414_));
 sky130_fd_sc_hd__a221o_1 _07977_ (.A1(_02410_),
    .A2(_02411_),
    .B1(_02412_),
    .B2(_02413_),
    .C1(_02414_),
    .X(_02415_));
 sky130_fd_sc_hd__o211a_1 _07978_ (.A1(_02405_),
    .A2(_02409_),
    .B1(_02415_),
    .C1(_02289_),
    .X(_02416_));
 sky130_fd_sc_hd__mux4_1 _07979_ (.A0(\regs[16][30] ),
    .A1(\regs[17][30] ),
    .A2(\regs[18][30] ),
    .A3(\regs[19][30] ),
    .S0(_02395_),
    .S1(_02351_),
    .X(_02417_));
 sky130_fd_sc_hd__buf_6 _07980_ (.A(_02329_),
    .X(_02418_));
 sky130_fd_sc_hd__mux4_1 _07981_ (.A0(\regs[20][30] ),
    .A1(\regs[21][30] ),
    .A2(\regs[22][30] ),
    .A3(\regs[23][30] ),
    .S0(_02348_),
    .S1(_02335_),
    .X(_02419_));
 sky130_fd_sc_hd__or2_1 _07982_ (.A(_02418_),
    .B(_02419_),
    .X(_02420_));
 sky130_fd_sc_hd__o211a_1 _07983_ (.A1(_02375_),
    .A2(_02417_),
    .B1(_02420_),
    .C1(_02361_),
    .X(_02421_));
 sky130_fd_sc_hd__buf_6 _07984_ (.A(_02408_),
    .X(_02422_));
 sky130_fd_sc_hd__buf_6 _07985_ (.A(_02367_),
    .X(_02423_));
 sky130_fd_sc_hd__mux4_1 _07986_ (.A0(\regs[12][30] ),
    .A1(\regs[13][30] ),
    .A2(\regs[14][30] ),
    .A3(\regs[15][30] ),
    .S0(_02303_),
    .S1(_02423_),
    .X(_02424_));
 sky130_fd_sc_hd__mux4_1 _07987_ (.A0(\regs[8][30] ),
    .A1(\regs[9][30] ),
    .A2(\regs[10][30] ),
    .A3(\regs[11][30] ),
    .S0(_02302_),
    .S1(_02367_),
    .X(_02425_));
 sky130_fd_sc_hd__or2_1 _07988_ (.A(_02293_),
    .B(_02425_),
    .X(_02426_));
 sky130_fd_sc_hd__o211a_1 _07989_ (.A1(_02422_),
    .A2(_02424_),
    .B1(_02426_),
    .C1(_02290_),
    .X(_02427_));
 sky130_fd_sc_hd__buf_8 _07990_ (.A(_02301_),
    .X(_02428_));
 sky130_fd_sc_hd__buf_6 _07991_ (.A(net9),
    .X(_02429_));
 sky130_fd_sc_hd__mux4_1 _07992_ (.A0(\regs[0][30] ),
    .A1(\regs[1][30] ),
    .A2(\regs[2][30] ),
    .A3(\regs[3][30] ),
    .S0(_02428_),
    .S1(_02429_),
    .X(_02430_));
 sky130_fd_sc_hd__mux4_1 _07993_ (.A0(\regs[4][30] ),
    .A1(\regs[5][30] ),
    .A2(\regs[6][30] ),
    .A3(\regs[7][30] ),
    .S0(_02332_),
    .S1(_02429_),
    .X(_02431_));
 sky130_fd_sc_hd__mux2_1 _07994_ (.A0(_02430_),
    .A1(_02431_),
    .S(_02414_),
    .X(_02432_));
 sky130_fd_sc_hd__buf_8 _07995_ (.A(net12),
    .X(_02433_));
 sky130_fd_sc_hd__a21o_1 _07996_ (.A1(_02362_),
    .A2(_02432_),
    .B1(_02433_),
    .X(_02434_));
 sky130_fd_sc_hd__o32a_1 _07997_ (.A1(_02286_),
    .A2(_02416_),
    .A3(_02421_),
    .B1(_02427_),
    .B2(_02434_),
    .X(_02435_));
 sky130_fd_sc_hd__mux2_1 _07998_ (.A0(\leorv32_alu.input1[30] ),
    .A1(_02435_),
    .S(_02324_),
    .X(_02436_));
 sky130_fd_sc_hd__clkbuf_1 _07999_ (.A(_02436_),
    .X(_01438_));
 sky130_fd_sc_hd__mux4_1 _08000_ (.A0(\regs[12][29] ),
    .A1(\regs[13][29] ),
    .A2(\regs[14][29] ),
    .A3(\regs[15][29] ),
    .S0(_02334_),
    .S1(_02337_),
    .X(_02437_));
 sky130_fd_sc_hd__or2_1 _08001_ (.A(_02331_),
    .B(_02437_),
    .X(_02438_));
 sky130_fd_sc_hd__mux4_2 _08002_ (.A0(\regs[8][29] ),
    .A1(\regs[9][29] ),
    .A2(\regs[10][29] ),
    .A3(\regs[11][29] ),
    .S0(_02341_),
    .S1(_02344_),
    .X(_02439_));
 sky130_fd_sc_hd__o21a_1 _08003_ (.A1(_02295_),
    .A2(_02439_),
    .B1(_02346_),
    .X(_02440_));
 sky130_fd_sc_hd__mux4_1 _08004_ (.A0(\regs[0][29] ),
    .A1(\regs[1][29] ),
    .A2(\regs[2][29] ),
    .A3(\regs[3][29] ),
    .S0(_02350_),
    .S1(_02352_),
    .X(_02441_));
 sky130_fd_sc_hd__mux4_1 _08005_ (.A0(\regs[4][29] ),
    .A1(\regs[5][29] ),
    .A2(\regs[6][29] ),
    .A3(\regs[7][29] ),
    .S0(_02355_),
    .S1(_02356_),
    .X(_02442_));
 sky130_fd_sc_hd__mux2_1 _08006_ (.A0(_02441_),
    .A1(_02442_),
    .S(_02359_),
    .X(_02443_));
 sky130_fd_sc_hd__a22o_1 _08007_ (.A1(_02438_),
    .A2(_02440_),
    .B1(_02443_),
    .B2(_02363_),
    .X(_02444_));
 sky130_fd_sc_hd__buf_6 _08008_ (.A(_02332_),
    .X(_02445_));
 sky130_fd_sc_hd__clkbuf_16 _08009_ (.A(_02445_),
    .X(_02446_));
 sky130_fd_sc_hd__buf_8 _08010_ (.A(_02343_),
    .X(_02447_));
 sky130_fd_sc_hd__mux4_1 _08011_ (.A0(\regs[20][29] ),
    .A1(\regs[21][29] ),
    .A2(\regs[22][29] ),
    .A3(\regs[23][29] ),
    .S0(_02446_),
    .S1(_02447_),
    .X(_02448_));
 sky130_fd_sc_hd__clkbuf_16 _08012_ (.A(_02333_),
    .X(_02449_));
 sky130_fd_sc_hd__buf_8 _08013_ (.A(_02343_),
    .X(_02450_));
 sky130_fd_sc_hd__mux4_1 _08014_ (.A0(\regs[16][29] ),
    .A1(\regs[17][29] ),
    .A2(\regs[18][29] ),
    .A3(\regs[19][29] ),
    .S0(_02449_),
    .S1(_02450_),
    .X(_02451_));
 sky130_fd_sc_hd__buf_8 _08015_ (.A(_02408_),
    .X(_02452_));
 sky130_fd_sc_hd__mux2_1 _08016_ (.A0(_02448_),
    .A1(_02451_),
    .S(_02452_),
    .X(_02453_));
 sky130_fd_sc_hd__buf_4 _08017_ (.A(_02336_),
    .X(_02454_));
 sky130_fd_sc_hd__clkbuf_8 _08018_ (.A(_02406_),
    .X(_02455_));
 sky130_fd_sc_hd__mux2_1 _08019_ (.A0(\regs[30][29] ),
    .A1(\regs[31][29] ),
    .S(_02455_),
    .X(_02456_));
 sky130_fd_sc_hd__and2_1 _08020_ (.A(_02454_),
    .B(_02456_),
    .X(_02457_));
 sky130_fd_sc_hd__buf_6 _08021_ (.A(_02301_),
    .X(_02458_));
 sky130_fd_sc_hd__buf_6 _08022_ (.A(_02458_),
    .X(_02459_));
 sky130_fd_sc_hd__mux2_1 _08023_ (.A0(\regs[28][29] ),
    .A1(\regs[29][29] ),
    .S(_02459_),
    .X(_02460_));
 sky130_fd_sc_hd__a21o_1 _08024_ (.A1(_02389_),
    .A2(_02460_),
    .B1(_02452_),
    .X(_02461_));
 sky130_fd_sc_hd__buf_8 _08025_ (.A(_02354_),
    .X(_02462_));
 sky130_fd_sc_hd__or2b_1 _08026_ (.A(\regs[27][29] ),
    .B_N(_02462_),
    .X(_02463_));
 sky130_fd_sc_hd__o21a_1 _08027_ (.A1(_02462_),
    .A2(\regs[26][29] ),
    .B1(_02368_),
    .X(_02464_));
 sky130_fd_sc_hd__mux2_1 _08028_ (.A0(\regs[24][29] ),
    .A1(\regs[25][29] ),
    .S(_02455_),
    .X(_02465_));
 sky130_fd_sc_hd__buf_4 _08029_ (.A(_02413_),
    .X(_02466_));
 sky130_fd_sc_hd__a221o_1 _08030_ (.A1(_02463_),
    .A2(_02464_),
    .B1(_02465_),
    .B2(_02466_),
    .C1(_02294_),
    .X(_02467_));
 sky130_fd_sc_hd__buf_4 _08031_ (.A(net11),
    .X(_02468_));
 sky130_fd_sc_hd__buf_6 _08032_ (.A(_02468_),
    .X(_02469_));
 sky130_fd_sc_hd__o211a_1 _08033_ (.A1(_02457_),
    .A2(_02461_),
    .B1(_02467_),
    .C1(_02469_),
    .X(_02470_));
 sky130_fd_sc_hd__buf_6 _08034_ (.A(_02399_),
    .X(_02471_));
 sky130_fd_sc_hd__a211o_1 _08035_ (.A1(_02366_),
    .A2(_02453_),
    .B1(_02470_),
    .C1(_02471_),
    .X(_02472_));
 sky130_fd_sc_hd__o221a_1 _08036_ (.A1(\leorv32_alu.input1[29] ),
    .A2(_02328_),
    .B1(_02288_),
    .B2(_02444_),
    .C1(_02472_),
    .X(_01437_));
 sky130_fd_sc_hd__mux2_1 _08037_ (.A0(\regs[30][28] ),
    .A1(\regs[31][28] ),
    .S(_02403_),
    .X(_02473_));
 sky130_fd_sc_hd__and2_1 _08038_ (.A(_02402_),
    .B(_02473_),
    .X(_02474_));
 sky130_fd_sc_hd__mux2_1 _08039_ (.A0(\regs[28][28] ),
    .A1(\regs[29][28] ),
    .S(_02406_),
    .X(_02475_));
 sky130_fd_sc_hd__a21o_1 _08040_ (.A1(_02413_),
    .A2(_02475_),
    .B1(_02408_),
    .X(_02476_));
 sky130_fd_sc_hd__or2b_1 _08041_ (.A(\regs[27][28] ),
    .B_N(_02380_),
    .X(_02477_));
 sky130_fd_sc_hd__o21a_1 _08042_ (.A1(_02380_),
    .A2(\regs[26][28] ),
    .B1(_02342_),
    .X(_02478_));
 sky130_fd_sc_hd__mux2_1 _08043_ (.A0(\regs[24][28] ),
    .A1(\regs[25][28] ),
    .S(_02302_),
    .X(_02479_));
 sky130_fd_sc_hd__a221o_1 _08044_ (.A1(_02477_),
    .A2(_02478_),
    .B1(_02479_),
    .B2(_02413_),
    .C1(_02414_),
    .X(_02480_));
 sky130_fd_sc_hd__o211a_1 _08045_ (.A1(_02474_),
    .A2(_02476_),
    .B1(_02480_),
    .C1(_02289_),
    .X(_02481_));
 sky130_fd_sc_hd__mux4_1 _08046_ (.A0(\regs[16][28] ),
    .A1(\regs[17][28] ),
    .A2(\regs[18][28] ),
    .A3(\regs[19][28] ),
    .S0(_02395_),
    .S1(_02351_),
    .X(_02482_));
 sky130_fd_sc_hd__mux4_1 _08047_ (.A0(\regs[20][28] ),
    .A1(\regs[21][28] ),
    .A2(\regs[22][28] ),
    .A3(\regs[23][28] ),
    .S0(_02348_),
    .S1(_02335_),
    .X(_02483_));
 sky130_fd_sc_hd__or2_1 _08048_ (.A(_02418_),
    .B(_02483_),
    .X(_02484_));
 sky130_fd_sc_hd__o211a_1 _08049_ (.A1(_02375_),
    .A2(_02482_),
    .B1(_02484_),
    .C1(_02361_),
    .X(_02485_));
 sky130_fd_sc_hd__mux4_1 _08050_ (.A0(\regs[12][28] ),
    .A1(\regs[13][28] ),
    .A2(\regs[14][28] ),
    .A3(\regs[15][28] ),
    .S0(_02303_),
    .S1(_02423_),
    .X(_02486_));
 sky130_fd_sc_hd__mux4_1 _08051_ (.A0(\regs[8][28] ),
    .A1(\regs[9][28] ),
    .A2(\regs[10][28] ),
    .A3(\regs[11][28] ),
    .S0(_02428_),
    .S1(_02367_),
    .X(_02487_));
 sky130_fd_sc_hd__or2_1 _08052_ (.A(_02293_),
    .B(_02487_),
    .X(_02488_));
 sky130_fd_sc_hd__o211a_1 _08053_ (.A1(_02422_),
    .A2(_02486_),
    .B1(_02488_),
    .C1(_02468_),
    .X(_02489_));
 sky130_fd_sc_hd__mux4_1 _08054_ (.A0(\regs[0][28] ),
    .A1(\regs[1][28] ),
    .A2(\regs[2][28] ),
    .A3(\regs[3][28] ),
    .S0(_02428_),
    .S1(_02429_),
    .X(_02490_));
 sky130_fd_sc_hd__mux4_1 _08055_ (.A0(\regs[4][28] ),
    .A1(\regs[5][28] ),
    .A2(\regs[6][28] ),
    .A3(\regs[7][28] ),
    .S0(_02332_),
    .S1(_02342_),
    .X(_02491_));
 sky130_fd_sc_hd__mux2_1 _08056_ (.A0(_02490_),
    .A1(_02491_),
    .S(_02414_),
    .X(_02492_));
 sky130_fd_sc_hd__a21o_1 _08057_ (.A1(_02362_),
    .A2(_02492_),
    .B1(_02433_),
    .X(_02493_));
 sky130_fd_sc_hd__o32a_2 _08058_ (.A1(_02286_),
    .A2(_02481_),
    .A3(_02485_),
    .B1(_02489_),
    .B2(_02493_),
    .X(_02494_));
 sky130_fd_sc_hd__mux2_1 _08059_ (.A0(_01736_),
    .A1(_02494_),
    .S(_02324_),
    .X(_02495_));
 sky130_fd_sc_hd__clkbuf_1 _08060_ (.A(_02495_),
    .X(_01436_));
 sky130_fd_sc_hd__mux4_1 _08061_ (.A0(\regs[12][27] ),
    .A1(\regs[13][27] ),
    .A2(\regs[14][27] ),
    .A3(\regs[15][27] ),
    .S0(_02334_),
    .S1(_02337_),
    .X(_02496_));
 sky130_fd_sc_hd__or2_1 _08062_ (.A(_02331_),
    .B(_02496_),
    .X(_02497_));
 sky130_fd_sc_hd__mux4_1 _08063_ (.A0(\regs[8][27] ),
    .A1(\regs[9][27] ),
    .A2(\regs[10][27] ),
    .A3(\regs[11][27] ),
    .S0(_02341_),
    .S1(_02344_),
    .X(_02498_));
 sky130_fd_sc_hd__o21a_1 _08064_ (.A1(_02295_),
    .A2(_02498_),
    .B1(_02346_),
    .X(_02499_));
 sky130_fd_sc_hd__mux4_1 _08065_ (.A0(\regs[0][27] ),
    .A1(\regs[1][27] ),
    .A2(\regs[2][27] ),
    .A3(\regs[3][27] ),
    .S0(_02350_),
    .S1(_02352_),
    .X(_02500_));
 sky130_fd_sc_hd__mux4_1 _08066_ (.A0(\regs[4][27] ),
    .A1(\regs[5][27] ),
    .A2(\regs[6][27] ),
    .A3(\regs[7][27] ),
    .S0(_02355_),
    .S1(_02356_),
    .X(_02501_));
 sky130_fd_sc_hd__mux2_1 _08067_ (.A0(_02500_),
    .A1(_02501_),
    .S(_02359_),
    .X(_02502_));
 sky130_fd_sc_hd__a22o_1 _08068_ (.A1(_02497_),
    .A2(_02499_),
    .B1(_02502_),
    .B2(_02363_),
    .X(_02503_));
 sky130_fd_sc_hd__mux4_1 _08069_ (.A0(\regs[16][27] ),
    .A1(\regs[17][27] ),
    .A2(\regs[18][27] ),
    .A3(\regs[19][27] ),
    .S0(_02304_),
    .S1(_02369_),
    .X(_02504_));
 sky130_fd_sc_hd__mux4_1 _08070_ (.A0(\regs[20][27] ),
    .A1(\regs[21][27] ),
    .A2(\regs[22][27] ),
    .A3(\regs[23][27] ),
    .S0(_02372_),
    .S1(_02373_),
    .X(_02505_));
 sky130_fd_sc_hd__mux2_1 _08071_ (.A0(_02504_),
    .A1(_02505_),
    .S(_02376_),
    .X(_02506_));
 sky130_fd_sc_hd__mux2_1 _08072_ (.A0(\regs[30][27] ),
    .A1(\regs[31][27] ),
    .S(_02392_),
    .X(_02507_));
 sky130_fd_sc_hd__clkbuf_8 _08073_ (.A(_02387_),
    .X(_02508_));
 sky130_fd_sc_hd__mux2_1 _08074_ (.A0(\regs[28][27] ),
    .A1(\regs[29][27] ),
    .S(_02333_),
    .X(_02509_));
 sky130_fd_sc_hd__a21o_1 _08075_ (.A1(_02508_),
    .A2(_02509_),
    .B1(_02330_),
    .X(_02510_));
 sky130_fd_sc_hd__a21o_1 _08076_ (.A1(_02299_),
    .A2(_02507_),
    .B1(_02510_),
    .X(_02511_));
 sky130_fd_sc_hd__or2b_1 _08077_ (.A(\regs[27][27] ),
    .B_N(_02381_),
    .X(_02512_));
 sky130_fd_sc_hd__o21a_1 _08078_ (.A1(_02381_),
    .A2(\regs[26][27] ),
    .B1(_02382_),
    .X(_02513_));
 sky130_fd_sc_hd__mux2_1 _08079_ (.A0(\regs[24][27] ),
    .A1(\regs[25][27] ),
    .S(_02459_),
    .X(_02514_));
 sky130_fd_sc_hd__clkbuf_8 _08080_ (.A(_02293_),
    .X(_02515_));
 sky130_fd_sc_hd__a221o_1 _08081_ (.A1(_02512_),
    .A2(_02513_),
    .B1(_02514_),
    .B2(_02466_),
    .C1(_02515_),
    .X(_02516_));
 sky130_fd_sc_hd__a31o_1 _08082_ (.A1(_02291_),
    .A2(_02511_),
    .A3(_02516_),
    .B1(_02399_),
    .X(_02517_));
 sky130_fd_sc_hd__a21o_1 _08083_ (.A1(_02366_),
    .A2(_02506_),
    .B1(_02517_),
    .X(_02518_));
 sky130_fd_sc_hd__o221a_1 _08084_ (.A1(\leorv32_alu.input1[27] ),
    .A2(_02328_),
    .B1(_02288_),
    .B2(_02503_),
    .C1(_02518_),
    .X(_01435_));
 sky130_fd_sc_hd__mux4_1 _08085_ (.A0(\regs[12][26] ),
    .A1(\regs[13][26] ),
    .A2(\regs[14][26] ),
    .A3(\regs[15][26] ),
    .S0(_02334_),
    .S1(_02337_),
    .X(_02519_));
 sky130_fd_sc_hd__or2_1 _08086_ (.A(_02331_),
    .B(_02519_),
    .X(_02520_));
 sky130_fd_sc_hd__mux4_1 _08087_ (.A0(\regs[8][26] ),
    .A1(\regs[9][26] ),
    .A2(\regs[10][26] ),
    .A3(\regs[11][26] ),
    .S0(_02341_),
    .S1(_02344_),
    .X(_02521_));
 sky130_fd_sc_hd__o21a_1 _08088_ (.A1(_02295_),
    .A2(_02521_),
    .B1(_02346_),
    .X(_02522_));
 sky130_fd_sc_hd__buf_8 _08089_ (.A(_02354_),
    .X(_02523_));
 sky130_fd_sc_hd__mux4_1 _08090_ (.A0(\regs[0][26] ),
    .A1(\regs[1][26] ),
    .A2(\regs[2][26] ),
    .A3(\regs[3][26] ),
    .S0(_02523_),
    .S1(_02352_),
    .X(_02524_));
 sky130_fd_sc_hd__mux4_1 _08091_ (.A0(\regs[4][26] ),
    .A1(\regs[5][26] ),
    .A2(\regs[6][26] ),
    .A3(\regs[7][26] ),
    .S0(_02355_),
    .S1(_02356_),
    .X(_02525_));
 sky130_fd_sc_hd__buf_6 _08092_ (.A(_02358_),
    .X(_02526_));
 sky130_fd_sc_hd__mux2_1 _08093_ (.A0(_02524_),
    .A1(_02525_),
    .S(_02526_),
    .X(_02527_));
 sky130_fd_sc_hd__a22o_1 _08094_ (.A1(_02520_),
    .A2(_02522_),
    .B1(_02527_),
    .B2(_02363_),
    .X(_02528_));
 sky130_fd_sc_hd__mux4_1 _08095_ (.A0(\regs[16][26] ),
    .A1(\regs[17][26] ),
    .A2(\regs[18][26] ),
    .A3(\regs[19][26] ),
    .S0(_02304_),
    .S1(_02369_),
    .X(_02529_));
 sky130_fd_sc_hd__mux4_1 _08096_ (.A0(\regs[20][26] ),
    .A1(\regs[21][26] ),
    .A2(\regs[22][26] ),
    .A3(\regs[23][26] ),
    .S0(_02372_),
    .S1(_02373_),
    .X(_02530_));
 sky130_fd_sc_hd__mux2_1 _08097_ (.A0(_02529_),
    .A1(_02530_),
    .S(_02376_),
    .X(_02531_));
 sky130_fd_sc_hd__or2b_1 _08098_ (.A(\regs[27][26] ),
    .B_N(_02378_),
    .X(_02532_));
 sky130_fd_sc_hd__o21a_1 _08099_ (.A1(_02381_),
    .A2(\regs[26][26] ),
    .B1(_02382_),
    .X(_02533_));
 sky130_fd_sc_hd__mux2_1 _08100_ (.A0(\regs[24][26] ),
    .A1(\regs[25][26] ),
    .S(_02384_),
    .X(_02534_));
 sky130_fd_sc_hd__a221o_1 _08101_ (.A1(_02532_),
    .A2(_02533_),
    .B1(_02534_),
    .B2(_02389_),
    .C1(_02390_),
    .X(_02535_));
 sky130_fd_sc_hd__mux2_1 _08102_ (.A0(\regs[30][26] ),
    .A1(\regs[31][26] ),
    .S(_02392_),
    .X(_02536_));
 sky130_fd_sc_hd__mux2_1 _08103_ (.A0(\regs[28][26] ),
    .A1(\regs[29][26] ),
    .S(_02395_),
    .X(_02537_));
 sky130_fd_sc_hd__buf_6 _08104_ (.A(_02329_),
    .X(_02538_));
 sky130_fd_sc_hd__a21o_1 _08105_ (.A1(_02394_),
    .A2(_02537_),
    .B1(_02538_),
    .X(_02539_));
 sky130_fd_sc_hd__a21o_1 _08106_ (.A1(_02299_),
    .A2(_02536_),
    .B1(_02539_),
    .X(_02540_));
 sky130_fd_sc_hd__a31o_1 _08107_ (.A1(_02291_),
    .A2(_02535_),
    .A3(_02540_),
    .B1(_02399_),
    .X(_02541_));
 sky130_fd_sc_hd__a21o_1 _08108_ (.A1(_02366_),
    .A2(_02531_),
    .B1(_02541_),
    .X(_02542_));
 sky130_fd_sc_hd__o221a_1 _08109_ (.A1(\leorv32_alu.input1[26] ),
    .A2(_02328_),
    .B1(_02288_),
    .B2(_02528_),
    .C1(_02542_),
    .X(_01434_));
 sky130_fd_sc_hd__buf_6 _08110_ (.A(_02251_),
    .X(_02543_));
 sky130_fd_sc_hd__mux4_1 _08111_ (.A0(\regs[12][25] ),
    .A1(\regs[13][25] ),
    .A2(\regs[14][25] ),
    .A3(\regs[15][25] ),
    .S0(_02340_),
    .S1(_02343_),
    .X(_02544_));
 sky130_fd_sc_hd__or2_1 _08112_ (.A(_02422_),
    .B(_02544_),
    .X(_02545_));
 sky130_fd_sc_hd__mux4_1 _08113_ (.A0(\regs[8][25] ),
    .A1(\regs[9][25] ),
    .A2(\regs[10][25] ),
    .A3(\regs[11][25] ),
    .S0(_02371_),
    .S1(_02402_),
    .X(_02546_));
 sky130_fd_sc_hd__o21a_1 _08114_ (.A1(_02515_),
    .A2(_02546_),
    .B1(_02468_),
    .X(_02547_));
 sky130_fd_sc_hd__mux4_1 _08115_ (.A0(\regs[0][25] ),
    .A1(\regs[1][25] ),
    .A2(\regs[2][25] ),
    .A3(\regs[3][25] ),
    .S0(_02340_),
    .S1(_02336_),
    .X(_02548_));
 sky130_fd_sc_hd__mux4_1 _08116_ (.A0(\regs[4][25] ),
    .A1(\regs[5][25] ),
    .A2(\regs[6][25] ),
    .A3(\regs[7][25] ),
    .S0(_02445_),
    .S1(_02336_),
    .X(_02549_));
 sky130_fd_sc_hd__buf_6 _08117_ (.A(_02414_),
    .X(_02550_));
 sky130_fd_sc_hd__mux2_1 _08118_ (.A0(_02548_),
    .A1(_02549_),
    .S(_02550_),
    .X(_02551_));
 sky130_fd_sc_hd__a22o_1 _08119_ (.A1(_02545_),
    .A2(_02547_),
    .B1(_02551_),
    .B2(_02365_),
    .X(_02552_));
 sky130_fd_sc_hd__buf_6 _08120_ (.A(_02302_),
    .X(_02553_));
 sky130_fd_sc_hd__mux4_1 _08121_ (.A0(\regs[16][25] ),
    .A1(\regs[17][25] ),
    .A2(\regs[18][25] ),
    .A3(\regs[19][25] ),
    .S0(_02553_),
    .S1(_02368_),
    .X(_02554_));
 sky130_fd_sc_hd__buf_6 _08122_ (.A(_02367_),
    .X(_02555_));
 sky130_fd_sc_hd__mux4_1 _08123_ (.A0(\regs[20][25] ),
    .A1(\regs[21][25] ),
    .A2(\regs[22][25] ),
    .A3(\regs[23][25] ),
    .S0(_02303_),
    .S1(_02555_),
    .X(_02556_));
 sky130_fd_sc_hd__mux2_1 _08124_ (.A0(_02554_),
    .A1(_02556_),
    .S(_02294_),
    .X(_02557_));
 sky130_fd_sc_hd__mux2_1 _08125_ (.A0(\regs[30][25] ),
    .A1(\regs[31][25] ),
    .S(_02349_),
    .X(_02558_));
 sky130_fd_sc_hd__mux2_1 _08126_ (.A0(\regs[28][25] ),
    .A1(\regs[29][25] ),
    .S(_02348_),
    .X(_02559_));
 sky130_fd_sc_hd__a21o_1 _08127_ (.A1(_02387_),
    .A2(_02559_),
    .B1(_02418_),
    .X(_02560_));
 sky130_fd_sc_hd__a21o_1 _08128_ (.A1(_02298_),
    .A2(_02558_),
    .B1(_02560_),
    .X(_02561_));
 sky130_fd_sc_hd__or2b_1 _08129_ (.A(\regs[27][25] ),
    .B_N(_02445_),
    .X(_02562_));
 sky130_fd_sc_hd__o21a_1 _08130_ (.A1(_02333_),
    .A2(\regs[26][25] ),
    .B1(_02297_),
    .X(_02563_));
 sky130_fd_sc_hd__mux2_1 _08131_ (.A0(\regs[24][25] ),
    .A1(\regs[25][25] ),
    .S(_02458_),
    .X(_02564_));
 sky130_fd_sc_hd__a221o_1 _08132_ (.A1(_02562_),
    .A2(_02563_),
    .B1(_02564_),
    .B2(_02388_),
    .C1(_02358_),
    .X(_02565_));
 sky130_fd_sc_hd__a31o_1 _08133_ (.A1(_02290_),
    .A2(_02561_),
    .A3(_02565_),
    .B1(_02286_),
    .X(_02566_));
 sky130_fd_sc_hd__a21o_1 _08134_ (.A1(_02365_),
    .A2(_02557_),
    .B1(_02566_),
    .X(_02567_));
 sky130_fd_sc_hd__o211a_2 _08135_ (.A1(_02433_),
    .A2(_02552_),
    .B1(_02567_),
    .C1(_02254_),
    .X(_02568_));
 sky130_fd_sc_hd__a21o_1 _08136_ (.A1(\leorv32_alu.input1[25] ),
    .A2(_02543_),
    .B1(_02568_),
    .X(_01433_));
 sky130_fd_sc_hd__buf_6 _08137_ (.A(_02362_),
    .X(_02569_));
 sky130_fd_sc_hd__mux4_1 _08138_ (.A0(\regs[4][24] ),
    .A1(\regs[5][24] ),
    .A2(\regs[6][24] ),
    .A3(\regs[7][24] ),
    .S0(_02462_),
    .S1(_02298_),
    .X(_02570_));
 sky130_fd_sc_hd__buf_8 _08139_ (.A(_02354_),
    .X(_02571_));
 sky130_fd_sc_hd__buf_8 _08140_ (.A(_02297_),
    .X(_02572_));
 sky130_fd_sc_hd__mux4_1 _08141_ (.A0(\regs[0][24] ),
    .A1(\regs[1][24] ),
    .A2(\regs[2][24] ),
    .A3(\regs[3][24] ),
    .S0(_02571_),
    .S1(_02572_),
    .X(_02573_));
 sky130_fd_sc_hd__mux2_1 _08142_ (.A0(_02570_),
    .A1(_02573_),
    .S(_02452_),
    .X(_02574_));
 sky130_fd_sc_hd__buf_8 _08143_ (.A(_02445_),
    .X(_02575_));
 sky130_fd_sc_hd__buf_6 _08144_ (.A(_02343_),
    .X(_02576_));
 sky130_fd_sc_hd__mux4_1 _08145_ (.A0(\regs[12][24] ),
    .A1(\regs[13][24] ),
    .A2(\regs[14][24] ),
    .A3(\regs[15][24] ),
    .S0(_02575_),
    .S1(_02576_),
    .X(_02577_));
 sky130_fd_sc_hd__or2_1 _08146_ (.A(_02331_),
    .B(_02577_),
    .X(_02578_));
 sky130_fd_sc_hd__mux4_1 _08147_ (.A0(\regs[8][24] ),
    .A1(\regs[9][24] ),
    .A2(\regs[10][24] ),
    .A3(\regs[11][24] ),
    .S0(_02372_),
    .S1(_02344_),
    .X(_02579_));
 sky130_fd_sc_hd__o21a_1 _08148_ (.A1(_02295_),
    .A2(_02579_),
    .B1(_02469_),
    .X(_02580_));
 sky130_fd_sc_hd__a22o_1 _08149_ (.A1(_02569_),
    .A2(_02574_),
    .B1(_02578_),
    .B2(_02580_),
    .X(_02581_));
 sky130_fd_sc_hd__buf_6 _08150_ (.A(_02362_),
    .X(_02582_));
 sky130_fd_sc_hd__mux4_1 _08151_ (.A0(\regs[16][24] ),
    .A1(\regs[17][24] ),
    .A2(\regs[18][24] ),
    .A3(\regs[19][24] ),
    .S0(_02446_),
    .S1(_02447_),
    .X(_02583_));
 sky130_fd_sc_hd__mux4_1 _08152_ (.A0(\regs[20][24] ),
    .A1(\regs[21][24] ),
    .A2(\regs[22][24] ),
    .A3(\regs[23][24] ),
    .S0(_02449_),
    .S1(_02450_),
    .X(_02584_));
 sky130_fd_sc_hd__mux2_1 _08153_ (.A0(_02583_),
    .A1(_02584_),
    .S(_02359_),
    .X(_02585_));
 sky130_fd_sc_hd__buf_4 _08154_ (.A(_02289_),
    .X(_02586_));
 sky130_fd_sc_hd__buf_6 _08155_ (.A(_02406_),
    .X(_02587_));
 sky130_fd_sc_hd__mux2_1 _08156_ (.A0(\regs[30][24] ),
    .A1(\regs[31][24] ),
    .S(_02587_),
    .X(_02588_));
 sky130_fd_sc_hd__mux2_1 _08157_ (.A0(\regs[28][24] ),
    .A1(\regs[29][24] ),
    .S(_02354_),
    .X(_02589_));
 sky130_fd_sc_hd__a21o_1 _08158_ (.A1(_02394_),
    .A2(_02589_),
    .B1(_02538_),
    .X(_02590_));
 sky130_fd_sc_hd__a21o_1 _08159_ (.A1(_02454_),
    .A2(_02588_),
    .B1(_02590_),
    .X(_02591_));
 sky130_fd_sc_hd__buf_6 _08160_ (.A(_02380_),
    .X(_02592_));
 sky130_fd_sc_hd__or2b_1 _08161_ (.A(\regs[27][24] ),
    .B_N(_02592_),
    .X(_02593_));
 sky130_fd_sc_hd__o21a_1 _08162_ (.A1(_02384_),
    .A2(\regs[26][24] ),
    .B1(_02555_),
    .X(_02594_));
 sky130_fd_sc_hd__mux2_1 _08163_ (.A0(\regs[24][24] ),
    .A1(\regs[25][24] ),
    .S(_02553_),
    .X(_02595_));
 sky130_fd_sc_hd__a221o_1 _08164_ (.A1(_02593_),
    .A2(_02594_),
    .B1(_02595_),
    .B2(_02508_),
    .C1(_02550_),
    .X(_02596_));
 sky130_fd_sc_hd__and3_1 _08165_ (.A(_02586_),
    .B(_02591_),
    .C(_02596_),
    .X(_02597_));
 sky130_fd_sc_hd__a211o_1 _08166_ (.A1(_02582_),
    .A2(_02585_),
    .B1(_02597_),
    .C1(_02471_),
    .X(_02598_));
 sky130_fd_sc_hd__o221a_1 _08167_ (.A1(\leorv32_alu.input1[24] ),
    .A2(_02328_),
    .B1(_02288_),
    .B2(_02581_),
    .C1(_02598_),
    .X(_01432_));
 sky130_fd_sc_hd__mux4_1 _08168_ (.A0(\regs[0][23] ),
    .A1(\regs[1][23] ),
    .A2(\regs[2][23] ),
    .A3(\regs[3][23] ),
    .S0(_02462_),
    .S1(_02298_),
    .X(_02599_));
 sky130_fd_sc_hd__mux4_1 _08169_ (.A0(\regs[4][23] ),
    .A1(\regs[5][23] ),
    .A2(\regs[6][23] ),
    .A3(\regs[7][23] ),
    .S0(_02571_),
    .S1(_02572_),
    .X(_02600_));
 sky130_fd_sc_hd__mux2_1 _08170_ (.A0(_02599_),
    .A1(_02600_),
    .S(_02390_),
    .X(_02601_));
 sky130_fd_sc_hd__mux4_1 _08171_ (.A0(\regs[12][23] ),
    .A1(\regs[13][23] ),
    .A2(\regs[14][23] ),
    .A3(\regs[15][23] ),
    .S0(_02575_),
    .S1(_02447_),
    .X(_02602_));
 sky130_fd_sc_hd__or2_1 _08172_ (.A(_02331_),
    .B(_02602_),
    .X(_02603_));
 sky130_fd_sc_hd__mux4_1 _08173_ (.A0(\regs[8][23] ),
    .A1(\regs[9][23] ),
    .A2(\regs[10][23] ),
    .A3(\regs[11][23] ),
    .S0(_02341_),
    .S1(_02344_),
    .X(_02604_));
 sky130_fd_sc_hd__o21a_1 _08174_ (.A1(_02295_),
    .A2(_02604_),
    .B1(_02469_),
    .X(_02605_));
 sky130_fd_sc_hd__a22o_1 _08175_ (.A1(_02569_),
    .A2(_02601_),
    .B1(_02603_),
    .B2(_02605_),
    .X(_02606_));
 sky130_fd_sc_hd__mux4_1 _08176_ (.A0(\regs[16][23] ),
    .A1(\regs[17][23] ),
    .A2(\regs[18][23] ),
    .A3(\regs[19][23] ),
    .S0(_02446_),
    .S1(_02447_),
    .X(_02607_));
 sky130_fd_sc_hd__mux4_1 _08177_ (.A0(\regs[20][23] ),
    .A1(\regs[21][23] ),
    .A2(\regs[22][23] ),
    .A3(\regs[23][23] ),
    .S0(_02449_),
    .S1(_02450_),
    .X(_02608_));
 sky130_fd_sc_hd__mux2_1 _08178_ (.A0(_02607_),
    .A1(_02608_),
    .S(_02359_),
    .X(_02609_));
 sky130_fd_sc_hd__mux2_1 _08179_ (.A0(\regs[30][23] ),
    .A1(\regs[31][23] ),
    .S(_02587_),
    .X(_02610_));
 sky130_fd_sc_hd__mux2_1 _08180_ (.A0(\regs[28][23] ),
    .A1(\regs[29][23] ),
    .S(_02354_),
    .X(_02611_));
 sky130_fd_sc_hd__a21o_1 _08181_ (.A1(_02394_),
    .A2(_02611_),
    .B1(_02538_),
    .X(_02612_));
 sky130_fd_sc_hd__a21o_1 _08182_ (.A1(_02454_),
    .A2(_02610_),
    .B1(_02612_),
    .X(_02613_));
 sky130_fd_sc_hd__or2b_1 _08183_ (.A(\regs[27][23] ),
    .B_N(_02592_),
    .X(_02614_));
 sky130_fd_sc_hd__o21a_1 _08184_ (.A1(_02384_),
    .A2(\regs[26][23] ),
    .B1(_02555_),
    .X(_02615_));
 sky130_fd_sc_hd__mux2_1 _08185_ (.A0(\regs[24][23] ),
    .A1(\regs[25][23] ),
    .S(_02553_),
    .X(_02616_));
 sky130_fd_sc_hd__a221o_1 _08186_ (.A1(_02614_),
    .A2(_02615_),
    .B1(_02616_),
    .B2(_02508_),
    .C1(_02550_),
    .X(_02617_));
 sky130_fd_sc_hd__and3_1 _08187_ (.A(_02586_),
    .B(_02613_),
    .C(_02617_),
    .X(_02618_));
 sky130_fd_sc_hd__a211o_1 _08188_ (.A1(_02582_),
    .A2(_02609_),
    .B1(_02618_),
    .C1(_02471_),
    .X(_02619_));
 sky130_fd_sc_hd__o221a_1 _08189_ (.A1(\leorv32_alu.input1[23] ),
    .A2(_02328_),
    .B1(_02288_),
    .B2(_02606_),
    .C1(_02619_),
    .X(_01431_));
 sky130_fd_sc_hd__clkbuf_4 _08190_ (.A(_02330_),
    .X(_02620_));
 sky130_fd_sc_hd__mux4_1 _08191_ (.A0(\regs[12][22] ),
    .A1(\regs[13][22] ),
    .A2(\regs[14][22] ),
    .A3(\regs[15][22] ),
    .S0(_02334_),
    .S1(_02337_),
    .X(_02621_));
 sky130_fd_sc_hd__or2_1 _08192_ (.A(_02620_),
    .B(_02621_),
    .X(_02622_));
 sky130_fd_sc_hd__buf_4 _08193_ (.A(_02294_),
    .X(_02623_));
 sky130_fd_sc_hd__mux4_1 _08194_ (.A0(\regs[8][22] ),
    .A1(\regs[9][22] ),
    .A2(\regs[10][22] ),
    .A3(\regs[11][22] ),
    .S0(_02341_),
    .S1(_02576_),
    .X(_02624_));
 sky130_fd_sc_hd__o21a_1 _08195_ (.A1(_02623_),
    .A2(_02624_),
    .B1(_02346_),
    .X(_02625_));
 sky130_fd_sc_hd__mux4_1 _08196_ (.A0(\regs[0][22] ),
    .A1(\regs[1][22] ),
    .A2(\regs[2][22] ),
    .A3(\regs[3][22] ),
    .S0(_02523_),
    .S1(_02352_),
    .X(_02626_));
 sky130_fd_sc_hd__mux4_1 _08197_ (.A0(\regs[4][22] ),
    .A1(\regs[5][22] ),
    .A2(\regs[6][22] ),
    .A3(\regs[7][22] ),
    .S0(_02355_),
    .S1(_02356_),
    .X(_02627_));
 sky130_fd_sc_hd__mux2_1 _08198_ (.A0(_02626_),
    .A1(_02627_),
    .S(_02526_),
    .X(_02628_));
 sky130_fd_sc_hd__a22o_1 _08199_ (.A1(_02622_),
    .A2(_02625_),
    .B1(_02628_),
    .B2(_02363_),
    .X(_02629_));
 sky130_fd_sc_hd__mux4_1 _08200_ (.A0(\regs[16][22] ),
    .A1(\regs[17][22] ),
    .A2(\regs[18][22] ),
    .A3(\regs[19][22] ),
    .S0(_02304_),
    .S1(_02369_),
    .X(_02630_));
 sky130_fd_sc_hd__mux4_1 _08201_ (.A0(\regs[20][22] ),
    .A1(\regs[21][22] ),
    .A2(\regs[22][22] ),
    .A3(\regs[23][22] ),
    .S0(_02372_),
    .S1(_02373_),
    .X(_02631_));
 sky130_fd_sc_hd__mux2_1 _08202_ (.A0(_02630_),
    .A1(_02631_),
    .S(_02376_),
    .X(_02632_));
 sky130_fd_sc_hd__or2b_1 _08203_ (.A(\regs[27][22] ),
    .B_N(_02378_),
    .X(_02633_));
 sky130_fd_sc_hd__o21a_1 _08204_ (.A1(_02381_),
    .A2(\regs[26][22] ),
    .B1(_02382_),
    .X(_02634_));
 sky130_fd_sc_hd__mux2_1 _08205_ (.A0(\regs[24][22] ),
    .A1(\regs[25][22] ),
    .S(_02459_),
    .X(_02635_));
 sky130_fd_sc_hd__a221o_1 _08206_ (.A1(_02633_),
    .A2(_02634_),
    .B1(_02635_),
    .B2(_02389_),
    .C1(_02515_),
    .X(_02636_));
 sky130_fd_sc_hd__mux2_1 _08207_ (.A0(\regs[30][22] ),
    .A1(\regs[31][22] ),
    .S(_02392_),
    .X(_02637_));
 sky130_fd_sc_hd__mux2_1 _08208_ (.A0(\regs[28][22] ),
    .A1(\regs[29][22] ),
    .S(_02395_),
    .X(_02638_));
 sky130_fd_sc_hd__a21o_1 _08209_ (.A1(_02394_),
    .A2(_02638_),
    .B1(_02538_),
    .X(_02639_));
 sky130_fd_sc_hd__a21o_1 _08210_ (.A1(_02299_),
    .A2(_02637_),
    .B1(_02639_),
    .X(_02640_));
 sky130_fd_sc_hd__a31o_1 _08211_ (.A1(_02291_),
    .A2(_02636_),
    .A3(_02640_),
    .B1(_02399_),
    .X(_02641_));
 sky130_fd_sc_hd__a21o_1 _08212_ (.A1(_02366_),
    .A2(_02632_),
    .B1(_02641_),
    .X(_02642_));
 sky130_fd_sc_hd__o221a_1 _08213_ (.A1(\leorv32_alu.input1[22] ),
    .A2(_02328_),
    .B1(_02288_),
    .B2(_02629_),
    .C1(_02642_),
    .X(_01430_));
 sky130_fd_sc_hd__buf_6 _08214_ (.A(_02351_),
    .X(_02643_));
 sky130_fd_sc_hd__mux4_1 _08215_ (.A0(\regs[12][21] ),
    .A1(\regs[13][21] ),
    .A2(\regs[14][21] ),
    .A3(\regs[15][21] ),
    .S0(_02334_),
    .S1(_02643_),
    .X(_02644_));
 sky130_fd_sc_hd__or2_1 _08216_ (.A(_02620_),
    .B(_02644_),
    .X(_02645_));
 sky130_fd_sc_hd__mux4_1 _08217_ (.A0(\regs[8][21] ),
    .A1(\regs[9][21] ),
    .A2(\regs[10][21] ),
    .A3(\regs[11][21] ),
    .S0(_02575_),
    .S1(_02576_),
    .X(_02646_));
 sky130_fd_sc_hd__o21a_1 _08218_ (.A1(_02623_),
    .A2(_02646_),
    .B1(_02346_),
    .X(_02647_));
 sky130_fd_sc_hd__mux4_1 _08219_ (.A0(\regs[0][21] ),
    .A1(\regs[1][21] ),
    .A2(\regs[2][21] ),
    .A3(\regs[3][21] ),
    .S0(_02523_),
    .S1(_02352_),
    .X(_02648_));
 sky130_fd_sc_hd__mux4_1 _08220_ (.A0(\regs[4][21] ),
    .A1(\regs[5][21] ),
    .A2(\regs[6][21] ),
    .A3(\regs[7][21] ),
    .S0(_02355_),
    .S1(_02356_),
    .X(_02649_));
 sky130_fd_sc_hd__mux2_1 _08221_ (.A0(_02648_),
    .A1(_02649_),
    .S(_02526_),
    .X(_02650_));
 sky130_fd_sc_hd__a22o_1 _08222_ (.A1(_02645_),
    .A2(_02647_),
    .B1(_02650_),
    .B2(_02363_),
    .X(_02651_));
 sky130_fd_sc_hd__mux4_1 _08223_ (.A0(\regs[20][21] ),
    .A1(\regs[21][21] ),
    .A2(\regs[22][21] ),
    .A3(\regs[23][21] ),
    .S0(_02446_),
    .S1(_02447_),
    .X(_02652_));
 sky130_fd_sc_hd__mux4_1 _08224_ (.A0(\regs[16][21] ),
    .A1(\regs[17][21] ),
    .A2(\regs[18][21] ),
    .A3(\regs[19][21] ),
    .S0(_02449_),
    .S1(_02450_),
    .X(_02653_));
 sky130_fd_sc_hd__mux2_1 _08225_ (.A0(_02652_),
    .A1(_02653_),
    .S(_02452_),
    .X(_02654_));
 sky130_fd_sc_hd__mux2_1 _08226_ (.A0(\regs[30][21] ),
    .A1(\regs[31][21] ),
    .S(_02455_),
    .X(_02655_));
 sky130_fd_sc_hd__and2_1 _08227_ (.A(_02454_),
    .B(_02655_),
    .X(_02656_));
 sky130_fd_sc_hd__mux2_1 _08228_ (.A0(\regs[28][21] ),
    .A1(\regs[29][21] ),
    .S(_02459_),
    .X(_02657_));
 sky130_fd_sc_hd__a21o_1 _08229_ (.A1(_02389_),
    .A2(_02657_),
    .B1(_02452_),
    .X(_02658_));
 sky130_fd_sc_hd__or2b_1 _08230_ (.A(\regs[27][21] ),
    .B_N(_02462_),
    .X(_02659_));
 sky130_fd_sc_hd__o21a_1 _08231_ (.A1(_02462_),
    .A2(\regs[26][21] ),
    .B1(_02368_),
    .X(_02660_));
 sky130_fd_sc_hd__mux2_1 _08232_ (.A0(\regs[24][21] ),
    .A1(\regs[25][21] ),
    .S(_02455_),
    .X(_02661_));
 sky130_fd_sc_hd__a221o_1 _08233_ (.A1(_02659_),
    .A2(_02660_),
    .B1(_02661_),
    .B2(_02466_),
    .C1(_02294_),
    .X(_02662_));
 sky130_fd_sc_hd__o211a_1 _08234_ (.A1(_02656_),
    .A2(_02658_),
    .B1(_02662_),
    .C1(_02469_),
    .X(_02663_));
 sky130_fd_sc_hd__a211o_1 _08235_ (.A1(_02582_),
    .A2(_02654_),
    .B1(_02663_),
    .C1(_02471_),
    .X(_02664_));
 sky130_fd_sc_hd__o221a_1 _08236_ (.A1(\leorv32_alu.input1[21] ),
    .A2(_02328_),
    .B1(_02288_),
    .B2(_02651_),
    .C1(_02664_),
    .X(_01429_));
 sky130_fd_sc_hd__mux2_1 _08237_ (.A0(\regs[30][20] ),
    .A1(\regs[31][20] ),
    .S(_02403_),
    .X(_02665_));
 sky130_fd_sc_hd__and2_1 _08238_ (.A(_02402_),
    .B(_02665_),
    .X(_02666_));
 sky130_fd_sc_hd__mux2_1 _08239_ (.A0(\regs[28][20] ),
    .A1(\regs[29][20] ),
    .S(_02403_),
    .X(_02667_));
 sky130_fd_sc_hd__a21o_1 _08240_ (.A1(_02413_),
    .A2(_02667_),
    .B1(_02408_),
    .X(_02668_));
 sky130_fd_sc_hd__or2b_1 _08241_ (.A(\regs[27][20] ),
    .B_N(_02380_),
    .X(_02669_));
 sky130_fd_sc_hd__o21a_1 _08242_ (.A1(_02406_),
    .A2(\regs[26][20] ),
    .B1(_02342_),
    .X(_02670_));
 sky130_fd_sc_hd__mux2_1 _08243_ (.A0(\regs[24][20] ),
    .A1(\regs[25][20] ),
    .S(_02302_),
    .X(_02671_));
 sky130_fd_sc_hd__a221o_1 _08244_ (.A1(_02669_),
    .A2(_02670_),
    .B1(_02671_),
    .B2(_02413_),
    .C1(_02414_),
    .X(_02672_));
 sky130_fd_sc_hd__o211a_1 _08245_ (.A1(_02666_),
    .A2(_02668_),
    .B1(_02672_),
    .C1(_02289_),
    .X(_02673_));
 sky130_fd_sc_hd__mux4_1 _08246_ (.A0(\regs[16][20] ),
    .A1(\regs[17][20] ),
    .A2(\regs[18][20] ),
    .A3(\regs[19][20] ),
    .S0(_02395_),
    .S1(_02351_),
    .X(_02674_));
 sky130_fd_sc_hd__mux4_1 _08247_ (.A0(\regs[20][20] ),
    .A1(\regs[21][20] ),
    .A2(\regs[22][20] ),
    .A3(\regs[23][20] ),
    .S0(_02348_),
    .S1(_02335_),
    .X(_02675_));
 sky130_fd_sc_hd__or2_1 _08248_ (.A(_02418_),
    .B(_02675_),
    .X(_02676_));
 sky130_fd_sc_hd__o211a_1 _08249_ (.A1(_02375_),
    .A2(_02674_),
    .B1(_02676_),
    .C1(_02361_),
    .X(_02677_));
 sky130_fd_sc_hd__mux4_1 _08250_ (.A0(\regs[12][20] ),
    .A1(\regs[13][20] ),
    .A2(\regs[14][20] ),
    .A3(\regs[15][20] ),
    .S0(_02303_),
    .S1(_02423_),
    .X(_02678_));
 sky130_fd_sc_hd__mux4_1 _08251_ (.A0(\regs[8][20] ),
    .A1(\regs[9][20] ),
    .A2(\regs[10][20] ),
    .A3(\regs[11][20] ),
    .S0(_02428_),
    .S1(_02367_),
    .X(_02679_));
 sky130_fd_sc_hd__or2_1 _08252_ (.A(_02293_),
    .B(_02679_),
    .X(_02680_));
 sky130_fd_sc_hd__o211a_1 _08253_ (.A1(_02422_),
    .A2(_02678_),
    .B1(_02680_),
    .C1(_02468_),
    .X(_02681_));
 sky130_fd_sc_hd__mux4_1 _08254_ (.A0(\regs[0][20] ),
    .A1(\regs[1][20] ),
    .A2(\regs[2][20] ),
    .A3(\regs[3][20] ),
    .S0(_02428_),
    .S1(_02429_),
    .X(_02682_));
 sky130_fd_sc_hd__mux4_1 _08255_ (.A0(\regs[4][20] ),
    .A1(\regs[5][20] ),
    .A2(\regs[6][20] ),
    .A3(\regs[7][20] ),
    .S0(_02332_),
    .S1(_02342_),
    .X(_02683_));
 sky130_fd_sc_hd__mux2_1 _08256_ (.A0(_02682_),
    .A1(_02683_),
    .S(_02414_),
    .X(_02684_));
 sky130_fd_sc_hd__a21o_1 _08257_ (.A1(_02362_),
    .A2(_02684_),
    .B1(_02433_),
    .X(_02685_));
 sky130_fd_sc_hd__o32a_2 _08258_ (.A1(_02286_),
    .A2(_02673_),
    .A3(_02677_),
    .B1(_02681_),
    .B2(_02685_),
    .X(_02686_));
 sky130_fd_sc_hd__mux2_1 _08259_ (.A0(\leorv32_alu.input1[20] ),
    .A1(_02686_),
    .S(_02324_),
    .X(_02687_));
 sky130_fd_sc_hd__clkbuf_1 _08260_ (.A(_02687_),
    .X(_01428_));
 sky130_fd_sc_hd__mux4_1 _08261_ (.A0(\regs[12][19] ),
    .A1(\regs[13][19] ),
    .A2(\regs[14][19] ),
    .A3(\regs[15][19] ),
    .S0(_02334_),
    .S1(_02643_),
    .X(_02688_));
 sky130_fd_sc_hd__or2_1 _08262_ (.A(_02620_),
    .B(_02688_),
    .X(_02689_));
 sky130_fd_sc_hd__mux4_2 _08263_ (.A0(\regs[8][19] ),
    .A1(\regs[9][19] ),
    .A2(\regs[10][19] ),
    .A3(\regs[11][19] ),
    .S0(_02575_),
    .S1(_02576_),
    .X(_02690_));
 sky130_fd_sc_hd__o21a_1 _08264_ (.A1(_02623_),
    .A2(_02690_),
    .B1(_02346_),
    .X(_02691_));
 sky130_fd_sc_hd__mux4_1 _08265_ (.A0(\regs[0][19] ),
    .A1(\regs[1][19] ),
    .A2(\regs[2][19] ),
    .A3(\regs[3][19] ),
    .S0(_02523_),
    .S1(_02352_),
    .X(_02692_));
 sky130_fd_sc_hd__mux4_1 _08266_ (.A0(\regs[4][19] ),
    .A1(\regs[5][19] ),
    .A2(\regs[6][19] ),
    .A3(\regs[7][19] ),
    .S0(_02355_),
    .S1(_02356_),
    .X(_02693_));
 sky130_fd_sc_hd__mux2_1 _08267_ (.A0(_02692_),
    .A1(_02693_),
    .S(_02526_),
    .X(_02694_));
 sky130_fd_sc_hd__a22o_2 _08268_ (.A1(_02689_),
    .A2(_02691_),
    .B1(_02694_),
    .B2(_02363_),
    .X(_02695_));
 sky130_fd_sc_hd__mux4_1 _08269_ (.A0(\regs[16][19] ),
    .A1(\regs[17][19] ),
    .A2(\regs[18][19] ),
    .A3(\regs[19][19] ),
    .S0(_02304_),
    .S1(_02369_),
    .X(_02696_));
 sky130_fd_sc_hd__mux4_1 _08270_ (.A0(\regs[20][19] ),
    .A1(\regs[21][19] ),
    .A2(\regs[22][19] ),
    .A3(\regs[23][19] ),
    .S0(_02372_),
    .S1(_02373_),
    .X(_02697_));
 sky130_fd_sc_hd__mux2_1 _08271_ (.A0(_02696_),
    .A1(_02697_),
    .S(_02376_),
    .X(_02698_));
 sky130_fd_sc_hd__mux2_1 _08272_ (.A0(\regs[30][19] ),
    .A1(\regs[31][19] ),
    .S(_02392_),
    .X(_02699_));
 sky130_fd_sc_hd__mux2_1 _08273_ (.A0(\regs[28][19] ),
    .A1(\regs[29][19] ),
    .S(_02333_),
    .X(_02700_));
 sky130_fd_sc_hd__a21o_1 _08274_ (.A1(_02508_),
    .A2(_02700_),
    .B1(_02330_),
    .X(_02701_));
 sky130_fd_sc_hd__a21o_1 _08275_ (.A1(_02299_),
    .A2(_02699_),
    .B1(_02701_),
    .X(_02702_));
 sky130_fd_sc_hd__or2b_1 _08276_ (.A(\regs[27][19] ),
    .B_N(_02381_),
    .X(_02703_));
 sky130_fd_sc_hd__o21a_1 _08277_ (.A1(_02334_),
    .A2(\regs[26][19] ),
    .B1(_02368_),
    .X(_02704_));
 sky130_fd_sc_hd__mux2_1 _08278_ (.A0(\regs[24][19] ),
    .A1(\regs[25][19] ),
    .S(_02459_),
    .X(_02705_));
 sky130_fd_sc_hd__a221o_1 _08279_ (.A1(_02703_),
    .A2(_02704_),
    .B1(_02705_),
    .B2(_02466_),
    .C1(_02515_),
    .X(_02706_));
 sky130_fd_sc_hd__a31o_1 _08280_ (.A1(_02291_),
    .A2(_02702_),
    .A3(_02706_),
    .B1(_02399_),
    .X(_02707_));
 sky130_fd_sc_hd__a21o_1 _08281_ (.A1(_02366_),
    .A2(_02698_),
    .B1(_02707_),
    .X(_02708_));
 sky130_fd_sc_hd__o221a_1 _08282_ (.A1(_01717_),
    .A2(_02328_),
    .B1(_02288_),
    .B2(_02695_),
    .C1(_02708_),
    .X(_01427_));
 sky130_fd_sc_hd__clkbuf_4 _08283_ (.A(_02287_),
    .X(_02709_));
 sky130_fd_sc_hd__mux4_1 _08284_ (.A0(\regs[12][18] ),
    .A1(\regs[13][18] ),
    .A2(\regs[14][18] ),
    .A3(\regs[15][18] ),
    .S0(_02334_),
    .S1(_02643_),
    .X(_02710_));
 sky130_fd_sc_hd__or2_1 _08285_ (.A(_02620_),
    .B(_02710_),
    .X(_02711_));
 sky130_fd_sc_hd__mux4_1 _08286_ (.A0(\regs[8][18] ),
    .A1(\regs[9][18] ),
    .A2(\regs[10][18] ),
    .A3(\regs[11][18] ),
    .S0(_02575_),
    .S1(_02576_),
    .X(_02712_));
 sky130_fd_sc_hd__o21a_1 _08287_ (.A1(_02623_),
    .A2(_02712_),
    .B1(_02346_),
    .X(_02713_));
 sky130_fd_sc_hd__mux4_1 _08288_ (.A0(\regs[0][18] ),
    .A1(\regs[1][18] ),
    .A2(\regs[2][18] ),
    .A3(\regs[3][18] ),
    .S0(_02523_),
    .S1(_02352_),
    .X(_02714_));
 sky130_fd_sc_hd__buf_4 _08289_ (.A(_02351_),
    .X(_02715_));
 sky130_fd_sc_hd__mux4_1 _08290_ (.A0(\regs[4][18] ),
    .A1(\regs[5][18] ),
    .A2(\regs[6][18] ),
    .A3(\regs[7][18] ),
    .S0(_02355_),
    .S1(_02715_),
    .X(_02716_));
 sky130_fd_sc_hd__mux2_1 _08291_ (.A0(_02714_),
    .A1(_02716_),
    .S(_02526_),
    .X(_02717_));
 sky130_fd_sc_hd__a22o_2 _08292_ (.A1(_02711_),
    .A2(_02713_),
    .B1(_02717_),
    .B2(_02363_),
    .X(_02718_));
 sky130_fd_sc_hd__mux4_1 _08293_ (.A0(\regs[16][18] ),
    .A1(\regs[17][18] ),
    .A2(\regs[18][18] ),
    .A3(\regs[19][18] ),
    .S0(_02304_),
    .S1(_02369_),
    .X(_02719_));
 sky130_fd_sc_hd__mux4_1 _08294_ (.A0(\regs[20][18] ),
    .A1(\regs[21][18] ),
    .A2(\regs[22][18] ),
    .A3(\regs[23][18] ),
    .S0(_02372_),
    .S1(_02373_),
    .X(_02720_));
 sky130_fd_sc_hd__mux2_1 _08295_ (.A0(_02719_),
    .A1(_02720_),
    .S(_02376_),
    .X(_02721_));
 sky130_fd_sc_hd__or2b_1 _08296_ (.A(\regs[27][18] ),
    .B_N(_02378_),
    .X(_02722_));
 sky130_fd_sc_hd__o21a_1 _08297_ (.A1(_02381_),
    .A2(\regs[26][18] ),
    .B1(_02382_),
    .X(_02723_));
 sky130_fd_sc_hd__mux2_1 _08298_ (.A0(\regs[24][18] ),
    .A1(\regs[25][18] ),
    .S(_02459_),
    .X(_02724_));
 sky130_fd_sc_hd__a221o_1 _08299_ (.A1(_02722_),
    .A2(_02723_),
    .B1(_02724_),
    .B2(_02389_),
    .C1(_02515_),
    .X(_02725_));
 sky130_fd_sc_hd__mux2_1 _08300_ (.A0(\regs[30][18] ),
    .A1(\regs[31][18] ),
    .S(_02392_),
    .X(_02726_));
 sky130_fd_sc_hd__mux2_1 _08301_ (.A0(\regs[28][18] ),
    .A1(\regs[29][18] ),
    .S(_02395_),
    .X(_02727_));
 sky130_fd_sc_hd__a21o_1 _08302_ (.A1(_02394_),
    .A2(_02727_),
    .B1(_02538_),
    .X(_02728_));
 sky130_fd_sc_hd__a21o_1 _08303_ (.A1(_02299_),
    .A2(_02726_),
    .B1(_02728_),
    .X(_02729_));
 sky130_fd_sc_hd__a31o_1 _08304_ (.A1(_02291_),
    .A2(_02725_),
    .A3(_02729_),
    .B1(_02399_),
    .X(_02730_));
 sky130_fd_sc_hd__a21o_1 _08305_ (.A1(_02366_),
    .A2(_02721_),
    .B1(_02730_),
    .X(_02731_));
 sky130_fd_sc_hd__o221a_1 _08306_ (.A1(_01867_),
    .A2(_02328_),
    .B1(_02709_),
    .B2(_02718_),
    .C1(_02731_),
    .X(_01426_));
 sky130_fd_sc_hd__mux4_1 _08307_ (.A0(\regs[12][17] ),
    .A1(\regs[13][17] ),
    .A2(\regs[14][17] ),
    .A3(\regs[15][17] ),
    .S0(_02340_),
    .S1(_02343_),
    .X(_02732_));
 sky130_fd_sc_hd__or2_1 _08308_ (.A(_02330_),
    .B(_02732_),
    .X(_02733_));
 sky130_fd_sc_hd__mux4_1 _08309_ (.A0(\regs[8][17] ),
    .A1(\regs[9][17] ),
    .A2(\regs[10][17] ),
    .A3(\regs[11][17] ),
    .S0(_02371_),
    .S1(_02402_),
    .X(_02734_));
 sky130_fd_sc_hd__o21a_1 _08310_ (.A1(_02515_),
    .A2(_02734_),
    .B1(_02468_),
    .X(_02735_));
 sky130_fd_sc_hd__mux4_1 _08311_ (.A0(\regs[0][17] ),
    .A1(\regs[1][17] ),
    .A2(\regs[2][17] ),
    .A3(\regs[3][17] ),
    .S0(_02340_),
    .S1(_02336_),
    .X(_02736_));
 sky130_fd_sc_hd__mux4_1 _08312_ (.A0(\regs[4][17] ),
    .A1(\regs[5][17] ),
    .A2(\regs[6][17] ),
    .A3(\regs[7][17] ),
    .S0(_02445_),
    .S1(_02336_),
    .X(_02737_));
 sky130_fd_sc_hd__mux2_1 _08313_ (.A0(_02736_),
    .A1(_02737_),
    .S(_02550_),
    .X(_02738_));
 sky130_fd_sc_hd__a22o_1 _08314_ (.A1(_02733_),
    .A2(_02735_),
    .B1(_02738_),
    .B2(_02365_),
    .X(_02739_));
 sky130_fd_sc_hd__mux4_1 _08315_ (.A0(\regs[16][17] ),
    .A1(\regs[17][17] ),
    .A2(\regs[18][17] ),
    .A3(\regs[19][17] ),
    .S0(_02553_),
    .S1(_02368_),
    .X(_02740_));
 sky130_fd_sc_hd__mux4_1 _08316_ (.A0(\regs[20][17] ),
    .A1(\regs[21][17] ),
    .A2(\regs[22][17] ),
    .A3(\regs[23][17] ),
    .S0(_02303_),
    .S1(_02555_),
    .X(_02741_));
 sky130_fd_sc_hd__mux2_1 _08317_ (.A0(_02740_),
    .A1(_02741_),
    .S(_02294_),
    .X(_02742_));
 sky130_fd_sc_hd__mux2_1 _08318_ (.A0(\regs[30][17] ),
    .A1(\regs[31][17] ),
    .S(_02349_),
    .X(_02743_));
 sky130_fd_sc_hd__mux2_1 _08319_ (.A0(\regs[28][17] ),
    .A1(\regs[29][17] ),
    .S(_02348_),
    .X(_02744_));
 sky130_fd_sc_hd__a21o_1 _08320_ (.A1(_02387_),
    .A2(_02744_),
    .B1(_02418_),
    .X(_02745_));
 sky130_fd_sc_hd__a21o_1 _08321_ (.A1(_02298_),
    .A2(_02743_),
    .B1(_02745_),
    .X(_02746_));
 sky130_fd_sc_hd__or2b_1 _08322_ (.A(\regs[27][17] ),
    .B_N(_02445_),
    .X(_02747_));
 sky130_fd_sc_hd__o21a_1 _08323_ (.A1(_02333_),
    .A2(\regs[26][17] ),
    .B1(_02367_),
    .X(_02748_));
 sky130_fd_sc_hd__mux2_1 _08324_ (.A0(\regs[24][17] ),
    .A1(\regs[25][17] ),
    .S(_02458_),
    .X(_02749_));
 sky130_fd_sc_hd__a221o_1 _08325_ (.A1(_02747_),
    .A2(_02748_),
    .B1(_02749_),
    .B2(_02388_),
    .C1(_02358_),
    .X(_02750_));
 sky130_fd_sc_hd__a31o_1 _08326_ (.A1(_02290_),
    .A2(_02746_),
    .A3(_02750_),
    .B1(_02285_),
    .X(_02751_));
 sky130_fd_sc_hd__a21o_1 _08327_ (.A1(_02365_),
    .A2(_02742_),
    .B1(_02751_),
    .X(_02752_));
 sky130_fd_sc_hd__o211a_1 _08328_ (.A1(_02433_),
    .A2(_02739_),
    .B1(_02752_),
    .C1(_02254_),
    .X(_02753_));
 sky130_fd_sc_hd__a21o_1 _08329_ (.A1(_01723_),
    .A2(_02543_),
    .B1(_02753_),
    .X(_01425_));
 sky130_fd_sc_hd__clkbuf_4 _08330_ (.A(_02255_),
    .X(_02754_));
 sky130_fd_sc_hd__mux4_1 _08331_ (.A0(\regs[12][16] ),
    .A1(\regs[13][16] ),
    .A2(\regs[14][16] ),
    .A3(\regs[15][16] ),
    .S0(_02350_),
    .S1(_02643_),
    .X(_02755_));
 sky130_fd_sc_hd__or2_1 _08332_ (.A(_02620_),
    .B(_02755_),
    .X(_02756_));
 sky130_fd_sc_hd__mux4_1 _08333_ (.A0(\regs[8][16] ),
    .A1(\regs[9][16] ),
    .A2(\regs[10][16] ),
    .A3(\regs[11][16] ),
    .S0(_02575_),
    .S1(_02576_),
    .X(_02757_));
 sky130_fd_sc_hd__o21a_1 _08334_ (.A1(_02623_),
    .A2(_02757_),
    .B1(_02586_),
    .X(_02758_));
 sky130_fd_sc_hd__mux4_1 _08335_ (.A0(\regs[0][16] ),
    .A1(\regs[1][16] ),
    .A2(\regs[2][16] ),
    .A3(\regs[3][16] ),
    .S0(_02523_),
    .S1(_02352_),
    .X(_02759_));
 sky130_fd_sc_hd__mux4_1 _08336_ (.A0(\regs[4][16] ),
    .A1(\regs[5][16] ),
    .A2(\regs[6][16] ),
    .A3(\regs[7][16] ),
    .S0(_02355_),
    .S1(_02715_),
    .X(_02760_));
 sky130_fd_sc_hd__mux2_1 _08337_ (.A0(_02759_),
    .A1(_02760_),
    .S(_02526_),
    .X(_02761_));
 sky130_fd_sc_hd__a22o_2 _08338_ (.A1(_02756_),
    .A2(_02758_),
    .B1(_02761_),
    .B2(_02363_),
    .X(_02762_));
 sky130_fd_sc_hd__mux4_1 _08339_ (.A0(\regs[20][16] ),
    .A1(\regs[21][16] ),
    .A2(\regs[22][16] ),
    .A3(\regs[23][16] ),
    .S0(_02446_),
    .S1(_02447_),
    .X(_02763_));
 sky130_fd_sc_hd__mux4_1 _08340_ (.A0(\regs[16][16] ),
    .A1(\regs[17][16] ),
    .A2(\regs[18][16] ),
    .A3(\regs[19][16] ),
    .S0(_02449_),
    .S1(_02450_),
    .X(_02764_));
 sky130_fd_sc_hd__mux2_1 _08341_ (.A0(_02763_),
    .A1(_02764_),
    .S(_02452_),
    .X(_02765_));
 sky130_fd_sc_hd__mux2_1 _08342_ (.A0(\regs[30][16] ),
    .A1(\regs[31][16] ),
    .S(_02455_),
    .X(_02766_));
 sky130_fd_sc_hd__and2_1 _08343_ (.A(_02454_),
    .B(_02766_),
    .X(_02767_));
 sky130_fd_sc_hd__mux2_1 _08344_ (.A0(\regs[28][16] ),
    .A1(\regs[29][16] ),
    .S(_02459_),
    .X(_02768_));
 sky130_fd_sc_hd__a21o_1 _08345_ (.A1(_02389_),
    .A2(_02768_),
    .B1(_02452_),
    .X(_02769_));
 sky130_fd_sc_hd__buf_4 _08346_ (.A(_02349_),
    .X(_02770_));
 sky130_fd_sc_hd__or2b_1 _08347_ (.A(\regs[27][16] ),
    .B_N(_02770_),
    .X(_02771_));
 sky130_fd_sc_hd__o21a_1 _08348_ (.A1(_02770_),
    .A2(\regs[26][16] ),
    .B1(_02368_),
    .X(_02772_));
 sky130_fd_sc_hd__mux2_1 _08349_ (.A0(\regs[24][16] ),
    .A1(\regs[25][16] ),
    .S(_02587_),
    .X(_02773_));
 sky130_fd_sc_hd__a221o_1 _08350_ (.A1(_02771_),
    .A2(_02772_),
    .B1(_02773_),
    .B2(_02466_),
    .C1(_02294_),
    .X(_02774_));
 sky130_fd_sc_hd__o211a_1 _08351_ (.A1(_02767_),
    .A2(_02769_),
    .B1(_02469_),
    .C1(_02774_),
    .X(_02775_));
 sky130_fd_sc_hd__a211o_1 _08352_ (.A1(_02582_),
    .A2(_02765_),
    .B1(_02775_),
    .C1(_02471_),
    .X(_02776_));
 sky130_fd_sc_hd__o221a_1 _08353_ (.A1(_01868_),
    .A2(_02754_),
    .B1(_02709_),
    .B2(_02762_),
    .C1(_02776_),
    .X(_01424_));
 sky130_fd_sc_hd__mux2_1 _08354_ (.A0(\regs[30][15] ),
    .A1(\regs[31][15] ),
    .S(_02403_),
    .X(_02777_));
 sky130_fd_sc_hd__and2_1 _08355_ (.A(_02402_),
    .B(_02777_),
    .X(_02778_));
 sky130_fd_sc_hd__mux2_1 _08356_ (.A0(\regs[28][15] ),
    .A1(\regs[29][15] ),
    .S(_02403_),
    .X(_02779_));
 sky130_fd_sc_hd__a21o_1 _08357_ (.A1(_02413_),
    .A2(_02779_),
    .B1(_02408_),
    .X(_02780_));
 sky130_fd_sc_hd__or2b_1 _08358_ (.A(\regs[27][15] ),
    .B_N(_02380_),
    .X(_02781_));
 sky130_fd_sc_hd__o21a_1 _08359_ (.A1(_02406_),
    .A2(\regs[26][15] ),
    .B1(_02342_),
    .X(_02782_));
 sky130_fd_sc_hd__mux2_1 _08360_ (.A0(\regs[24][15] ),
    .A1(\regs[25][15] ),
    .S(_02302_),
    .X(_02783_));
 sky130_fd_sc_hd__a221o_1 _08361_ (.A1(_02781_),
    .A2(_02782_),
    .B1(_02783_),
    .B2(_02413_),
    .C1(net10),
    .X(_02784_));
 sky130_fd_sc_hd__o211a_1 _08362_ (.A1(_02778_),
    .A2(_02780_),
    .B1(_02784_),
    .C1(_02289_),
    .X(_02785_));
 sky130_fd_sc_hd__mux4_1 _08363_ (.A0(\regs[16][15] ),
    .A1(\regs[17][15] ),
    .A2(\regs[18][15] ),
    .A3(\regs[19][15] ),
    .S0(_02349_),
    .S1(_02351_),
    .X(_02786_));
 sky130_fd_sc_hd__mux4_1 _08364_ (.A0(\regs[20][15] ),
    .A1(\regs[21][15] ),
    .A2(\regs[22][15] ),
    .A3(\regs[23][15] ),
    .S0(_02348_),
    .S1(_02335_),
    .X(_02787_));
 sky130_fd_sc_hd__or2_1 _08365_ (.A(_02418_),
    .B(_02787_),
    .X(_02788_));
 sky130_fd_sc_hd__o211a_1 _08366_ (.A1(_02375_),
    .A2(_02786_),
    .B1(_02788_),
    .C1(_02361_),
    .X(_02789_));
 sky130_fd_sc_hd__mux4_1 _08367_ (.A0(\regs[12][15] ),
    .A1(\regs[13][15] ),
    .A2(\regs[14][15] ),
    .A3(\regs[15][15] ),
    .S0(_02371_),
    .S1(_02423_),
    .X(_02790_));
 sky130_fd_sc_hd__mux4_1 _08368_ (.A0(\regs[8][15] ),
    .A1(\regs[9][15] ),
    .A2(\regs[10][15] ),
    .A3(\regs[11][15] ),
    .S0(_02428_),
    .S1(_02429_),
    .X(_02791_));
 sky130_fd_sc_hd__or2_1 _08369_ (.A(_02293_),
    .B(_02791_),
    .X(_02792_));
 sky130_fd_sc_hd__o211a_1 _08370_ (.A1(_02422_),
    .A2(_02790_),
    .B1(_02792_),
    .C1(_02468_),
    .X(_02793_));
 sky130_fd_sc_hd__mux4_1 _08371_ (.A0(\regs[0][15] ),
    .A1(\regs[1][15] ),
    .A2(\regs[2][15] ),
    .A3(\regs[3][15] ),
    .S0(_02428_),
    .S1(_02429_),
    .X(_02794_));
 sky130_fd_sc_hd__mux4_1 _08372_ (.A0(\regs[4][15] ),
    .A1(\regs[5][15] ),
    .A2(\regs[6][15] ),
    .A3(\regs[7][15] ),
    .S0(_02332_),
    .S1(_02342_),
    .X(_02795_));
 sky130_fd_sc_hd__mux2_1 _08373_ (.A0(_02794_),
    .A1(_02795_),
    .S(_02414_),
    .X(_02796_));
 sky130_fd_sc_hd__a21o_1 _08374_ (.A1(_02362_),
    .A2(_02796_),
    .B1(net12),
    .X(_02797_));
 sky130_fd_sc_hd__o32a_1 _08375_ (.A1(_02286_),
    .A2(_02785_),
    .A3(_02789_),
    .B1(_02793_),
    .B2(_02797_),
    .X(_02798_));
 sky130_fd_sc_hd__mux2_1 _08376_ (.A0(_01870_),
    .A1(_02798_),
    .S(_02324_),
    .X(_02799_));
 sky130_fd_sc_hd__clkbuf_1 _08377_ (.A(_02799_),
    .X(_01423_));
 sky130_fd_sc_hd__mux4_1 _08378_ (.A0(\regs[12][14] ),
    .A1(\regs[13][14] ),
    .A2(\regs[14][14] ),
    .A3(\regs[15][14] ),
    .S0(_02350_),
    .S1(_02643_),
    .X(_02800_));
 sky130_fd_sc_hd__or2_1 _08379_ (.A(_02620_),
    .B(_02800_),
    .X(_02801_));
 sky130_fd_sc_hd__mux4_1 _08380_ (.A0(\regs[8][14] ),
    .A1(\regs[9][14] ),
    .A2(\regs[10][14] ),
    .A3(\regs[11][14] ),
    .S0(_02575_),
    .S1(_02576_),
    .X(_02802_));
 sky130_fd_sc_hd__o21a_1 _08381_ (.A1(_02623_),
    .A2(_02802_),
    .B1(_02586_),
    .X(_02803_));
 sky130_fd_sc_hd__mux4_1 _08382_ (.A0(\regs[0][14] ),
    .A1(\regs[1][14] ),
    .A2(\regs[2][14] ),
    .A3(\regs[3][14] ),
    .S0(_02523_),
    .S1(_02352_),
    .X(_02804_));
 sky130_fd_sc_hd__mux4_1 _08383_ (.A0(\regs[4][14] ),
    .A1(\regs[5][14] ),
    .A2(\regs[6][14] ),
    .A3(\regs[7][14] ),
    .S0(_02355_),
    .S1(_02715_),
    .X(_02805_));
 sky130_fd_sc_hd__mux2_1 _08384_ (.A0(_02804_),
    .A1(_02805_),
    .S(_02526_),
    .X(_02806_));
 sky130_fd_sc_hd__a22o_2 _08385_ (.A1(_02801_),
    .A2(_02803_),
    .B1(_02806_),
    .B2(_02569_),
    .X(_02807_));
 sky130_fd_sc_hd__mux4_1 _08386_ (.A0(\regs[16][14] ),
    .A1(\regs[17][14] ),
    .A2(\regs[18][14] ),
    .A3(\regs[19][14] ),
    .S0(_02304_),
    .S1(_02369_),
    .X(_02808_));
 sky130_fd_sc_hd__mux4_1 _08387_ (.A0(\regs[20][14] ),
    .A1(\regs[21][14] ),
    .A2(\regs[22][14] ),
    .A3(\regs[23][14] ),
    .S0(_02372_),
    .S1(_02373_),
    .X(_02809_));
 sky130_fd_sc_hd__mux2_1 _08388_ (.A0(_02808_),
    .A1(_02809_),
    .S(_02376_),
    .X(_02810_));
 sky130_fd_sc_hd__mux2_1 _08389_ (.A0(\regs[30][14] ),
    .A1(\regs[31][14] ),
    .S(_02392_),
    .X(_02811_));
 sky130_fd_sc_hd__mux2_1 _08390_ (.A0(\regs[28][14] ),
    .A1(\regs[29][14] ),
    .S(_02395_),
    .X(_02812_));
 sky130_fd_sc_hd__a21o_1 _08391_ (.A1(_02508_),
    .A2(_02812_),
    .B1(_02330_),
    .X(_02813_));
 sky130_fd_sc_hd__a21o_1 _08392_ (.A1(_02299_),
    .A2(_02811_),
    .B1(_02813_),
    .X(_02814_));
 sky130_fd_sc_hd__or2b_1 _08393_ (.A(\regs[27][14] ),
    .B_N(_02381_),
    .X(_02815_));
 sky130_fd_sc_hd__o21a_1 _08394_ (.A1(_02334_),
    .A2(\regs[26][14] ),
    .B1(_02368_),
    .X(_02816_));
 sky130_fd_sc_hd__mux2_1 _08395_ (.A0(\regs[24][14] ),
    .A1(\regs[25][14] ),
    .S(_02459_),
    .X(_02817_));
 sky130_fd_sc_hd__a221o_1 _08396_ (.A1(_02815_),
    .A2(_02816_),
    .B1(_02817_),
    .B2(_02466_),
    .C1(_02515_),
    .X(_02818_));
 sky130_fd_sc_hd__a31o_1 _08397_ (.A1(_02291_),
    .A2(_02814_),
    .A3(_02818_),
    .B1(_02399_),
    .X(_02819_));
 sky130_fd_sc_hd__a21o_1 _08398_ (.A1(_02366_),
    .A2(_02810_),
    .B1(_02819_),
    .X(_02820_));
 sky130_fd_sc_hd__o221a_1 _08399_ (.A1(_01871_),
    .A2(_02754_),
    .B1(_02709_),
    .B2(_02807_),
    .C1(_02820_),
    .X(_01422_));
 sky130_fd_sc_hd__mux4_1 _08400_ (.A0(\regs[12][13] ),
    .A1(\regs[13][13] ),
    .A2(\regs[14][13] ),
    .A3(\regs[15][13] ),
    .S0(_02350_),
    .S1(_02643_),
    .X(_02821_));
 sky130_fd_sc_hd__or2_1 _08401_ (.A(_02620_),
    .B(_02821_),
    .X(_02822_));
 sky130_fd_sc_hd__mux4_1 _08402_ (.A0(\regs[8][13] ),
    .A1(\regs[9][13] ),
    .A2(\regs[10][13] ),
    .A3(\regs[11][13] ),
    .S0(_02575_),
    .S1(_02576_),
    .X(_02823_));
 sky130_fd_sc_hd__o21a_1 _08403_ (.A1(_02623_),
    .A2(_02823_),
    .B1(_02586_),
    .X(_02824_));
 sky130_fd_sc_hd__mux4_1 _08404_ (.A0(\regs[0][13] ),
    .A1(\regs[1][13] ),
    .A2(\regs[2][13] ),
    .A3(\regs[3][13] ),
    .S0(_02523_),
    .S1(_02356_),
    .X(_02825_));
 sky130_fd_sc_hd__mux4_1 _08405_ (.A0(\regs[4][13] ),
    .A1(\regs[5][13] ),
    .A2(\regs[6][13] ),
    .A3(\regs[7][13] ),
    .S0(_02392_),
    .S1(_02715_),
    .X(_02826_));
 sky130_fd_sc_hd__mux2_1 _08406_ (.A0(_02825_),
    .A1(_02826_),
    .S(_02526_),
    .X(_02827_));
 sky130_fd_sc_hd__a22o_2 _08407_ (.A1(_02822_),
    .A2(_02824_),
    .B1(_02827_),
    .B2(_02569_),
    .X(_02828_));
 sky130_fd_sc_hd__mux4_1 _08408_ (.A0(\regs[16][13] ),
    .A1(\regs[17][13] ),
    .A2(\regs[18][13] ),
    .A3(\regs[19][13] ),
    .S0(_02304_),
    .S1(_02369_),
    .X(_02829_));
 sky130_fd_sc_hd__mux4_1 _08409_ (.A0(\regs[20][13] ),
    .A1(\regs[21][13] ),
    .A2(\regs[22][13] ),
    .A3(\regs[23][13] ),
    .S0(_02372_),
    .S1(_02373_),
    .X(_02830_));
 sky130_fd_sc_hd__mux2_1 _08410_ (.A0(_02829_),
    .A1(_02830_),
    .S(_02376_),
    .X(_02831_));
 sky130_fd_sc_hd__or2b_1 _08411_ (.A(\regs[27][13] ),
    .B_N(_02378_),
    .X(_02832_));
 sky130_fd_sc_hd__o21a_1 _08412_ (.A1(_02381_),
    .A2(\regs[26][13] ),
    .B1(_02382_),
    .X(_02833_));
 sky130_fd_sc_hd__mux2_1 _08413_ (.A0(\regs[24][13] ),
    .A1(\regs[25][13] ),
    .S(_02459_),
    .X(_02834_));
 sky130_fd_sc_hd__a221o_1 _08414_ (.A1(_02832_),
    .A2(_02833_),
    .B1(_02834_),
    .B2(_02389_),
    .C1(_02515_),
    .X(_02835_));
 sky130_fd_sc_hd__mux2_1 _08415_ (.A0(\regs[30][13] ),
    .A1(\regs[31][13] ),
    .S(_02770_),
    .X(_02836_));
 sky130_fd_sc_hd__mux2_1 _08416_ (.A0(\regs[28][13] ),
    .A1(\regs[29][13] ),
    .S(_02395_),
    .X(_02837_));
 sky130_fd_sc_hd__a21o_1 _08417_ (.A1(_02394_),
    .A2(_02837_),
    .B1(_02538_),
    .X(_02838_));
 sky130_fd_sc_hd__a21o_1 _08418_ (.A1(_02299_),
    .A2(_02836_),
    .B1(_02838_),
    .X(_02839_));
 sky130_fd_sc_hd__a31o_1 _08419_ (.A1(_02291_),
    .A2(_02835_),
    .A3(_02839_),
    .B1(_02399_),
    .X(_02840_));
 sky130_fd_sc_hd__a21o_1 _08420_ (.A1(_02366_),
    .A2(_02831_),
    .B1(_02840_),
    .X(_02841_));
 sky130_fd_sc_hd__o221a_1 _08421_ (.A1(_01872_),
    .A2(_02754_),
    .B1(_02709_),
    .B2(_02828_),
    .C1(_02841_),
    .X(_01421_));
 sky130_fd_sc_hd__mux4_1 _08422_ (.A0(\regs[16][12] ),
    .A1(\regs[17][12] ),
    .A2(\regs[18][12] ),
    .A3(\regs[19][12] ),
    .S0(_02770_),
    .S1(_02715_),
    .X(_02842_));
 sky130_fd_sc_hd__mux4_1 _08423_ (.A0(\regs[20][12] ),
    .A1(\regs[21][12] ),
    .A2(\regs[22][12] ),
    .A3(\regs[23][12] ),
    .S0(_02770_),
    .S1(_02715_),
    .X(_02843_));
 sky130_fd_sc_hd__mux2_1 _08424_ (.A0(_02842_),
    .A1(_02843_),
    .S(_02390_),
    .X(_02844_));
 sky130_fd_sc_hd__mux2_1 _08425_ (.A0(\regs[30][12] ),
    .A1(\regs[31][12] ),
    .S(_02455_),
    .X(_02845_));
 sky130_fd_sc_hd__and2_1 _08426_ (.A(_02369_),
    .B(_02845_),
    .X(_02846_));
 sky130_fd_sc_hd__mux2_1 _08427_ (.A0(\regs[28][12] ),
    .A1(\regs[29][12] ),
    .S(_02455_),
    .X(_02847_));
 sky130_fd_sc_hd__a21o_1 _08428_ (.A1(_02466_),
    .A2(_02847_),
    .B1(_02422_),
    .X(_02848_));
 sky130_fd_sc_hd__or2b_1 _08429_ (.A(\regs[27][12] ),
    .B_N(_02592_),
    .X(_02849_));
 sky130_fd_sc_hd__o21a_1 _08430_ (.A1(_02592_),
    .A2(\regs[26][12] ),
    .B1(_02555_),
    .X(_02850_));
 sky130_fd_sc_hd__mux2_1 _08431_ (.A0(\regs[24][12] ),
    .A1(\regs[25][12] ),
    .S(_02553_),
    .X(_02851_));
 sky130_fd_sc_hd__a221o_1 _08432_ (.A1(_02849_),
    .A2(_02850_),
    .B1(_02851_),
    .B2(_02466_),
    .C1(_02375_),
    .X(_02852_));
 sky130_fd_sc_hd__o211a_1 _08433_ (.A1(_02846_),
    .A2(_02848_),
    .B1(_02852_),
    .C1(_02346_),
    .X(_02853_));
 sky130_fd_sc_hd__a211o_1 _08434_ (.A1(_02582_),
    .A2(_02844_),
    .B1(_02853_),
    .C1(_02286_),
    .X(_02854_));
 sky130_fd_sc_hd__mux4_1 _08435_ (.A0(\regs[12][12] ),
    .A1(\regs[13][12] ),
    .A2(\regs[14][12] ),
    .A3(\regs[15][12] ),
    .S0(_02462_),
    .S1(_02298_),
    .X(_02855_));
 sky130_fd_sc_hd__or2_1 _08436_ (.A(_02620_),
    .B(_02855_),
    .X(_02856_));
 sky130_fd_sc_hd__mux4_1 _08437_ (.A0(\regs[8][12] ),
    .A1(\regs[9][12] ),
    .A2(\regs[10][12] ),
    .A3(\regs[11][12] ),
    .S0(_02350_),
    .S1(_02643_),
    .X(_02857_));
 sky130_fd_sc_hd__o21a_1 _08438_ (.A1(_02376_),
    .A2(_02857_),
    .B1(_02290_),
    .X(_02858_));
 sky130_fd_sc_hd__mux4_1 _08439_ (.A0(\regs[0][12] ),
    .A1(\regs[1][12] ),
    .A2(\regs[2][12] ),
    .A3(\regs[3][12] ),
    .S0(_02571_),
    .S1(_02572_),
    .X(_02859_));
 sky130_fd_sc_hd__mux4_1 _08440_ (.A0(\regs[4][12] ),
    .A1(\regs[5][12] ),
    .A2(\regs[6][12] ),
    .A3(\regs[7][12] ),
    .S0(_02592_),
    .S1(_02382_),
    .X(_02860_));
 sky130_fd_sc_hd__mux2_1 _08441_ (.A0(_02859_),
    .A1(_02860_),
    .S(_02390_),
    .X(_02861_));
 sky130_fd_sc_hd__a221o_2 _08442_ (.A1(_02856_),
    .A2(_02858_),
    .B1(_02861_),
    .B2(_02365_),
    .C1(_02433_),
    .X(_02862_));
 sky130_fd_sc_hd__and2_1 _08443_ (.A(_01747_),
    .B(_02543_),
    .X(_02863_));
 sky130_fd_sc_hd__a31o_1 _08444_ (.A1(_00001_),
    .A2(_02854_),
    .A3(_02862_),
    .B1(_02863_),
    .X(_01420_));
 sky130_fd_sc_hd__mux4_1 _08445_ (.A0(\regs[12][11] ),
    .A1(\regs[13][11] ),
    .A2(\regs[14][11] ),
    .A3(\regs[15][11] ),
    .S0(_02350_),
    .S1(_02643_),
    .X(_02864_));
 sky130_fd_sc_hd__or2_1 _08446_ (.A(_02620_),
    .B(_02864_),
    .X(_02865_));
 sky130_fd_sc_hd__mux4_1 _08447_ (.A0(\regs[8][11] ),
    .A1(\regs[9][11] ),
    .A2(\regs[10][11] ),
    .A3(\regs[11][11] ),
    .S0(_02575_),
    .S1(_02576_),
    .X(_02866_));
 sky130_fd_sc_hd__o21a_1 _08448_ (.A1(_02623_),
    .A2(_02866_),
    .B1(_02586_),
    .X(_02867_));
 sky130_fd_sc_hd__mux4_1 _08449_ (.A0(\regs[0][11] ),
    .A1(\regs[1][11] ),
    .A2(\regs[2][11] ),
    .A3(\regs[3][11] ),
    .S0(_02523_),
    .S1(_02356_),
    .X(_02868_));
 sky130_fd_sc_hd__mux4_1 _08450_ (.A0(\regs[4][11] ),
    .A1(\regs[5][11] ),
    .A2(\regs[6][11] ),
    .A3(\regs[7][11] ),
    .S0(_02392_),
    .S1(_02715_),
    .X(_02869_));
 sky130_fd_sc_hd__mux2_1 _08451_ (.A0(_02868_),
    .A1(_02869_),
    .S(_02526_),
    .X(_02870_));
 sky130_fd_sc_hd__a22o_2 _08452_ (.A1(_02865_),
    .A2(_02867_),
    .B1(_02870_),
    .B2(_02569_),
    .X(_02871_));
 sky130_fd_sc_hd__mux4_1 _08453_ (.A0(\regs[16][11] ),
    .A1(\regs[17][11] ),
    .A2(\regs[18][11] ),
    .A3(\regs[19][11] ),
    .S0(_02304_),
    .S1(_02373_),
    .X(_02872_));
 sky130_fd_sc_hd__mux4_1 _08454_ (.A0(\regs[20][11] ),
    .A1(\regs[21][11] ),
    .A2(\regs[22][11] ),
    .A3(\regs[23][11] ),
    .S0(_02372_),
    .S1(_02373_),
    .X(_02873_));
 sky130_fd_sc_hd__mux2_1 _08455_ (.A0(_02872_),
    .A1(_02873_),
    .S(_02376_),
    .X(_02874_));
 sky130_fd_sc_hd__or2b_1 _08456_ (.A(\regs[27][11] ),
    .B_N(_02378_),
    .X(_02875_));
 sky130_fd_sc_hd__o21a_1 _08457_ (.A1(_02381_),
    .A2(\regs[26][11] ),
    .B1(_02382_),
    .X(_02876_));
 sky130_fd_sc_hd__mux2_1 _08458_ (.A0(\regs[24][11] ),
    .A1(\regs[25][11] ),
    .S(_02459_),
    .X(_02877_));
 sky130_fd_sc_hd__a221o_1 _08459_ (.A1(_02875_),
    .A2(_02876_),
    .B1(_02877_),
    .B2(_02389_),
    .C1(_02515_),
    .X(_02878_));
 sky130_fd_sc_hd__mux2_1 _08460_ (.A0(\regs[30][11] ),
    .A1(\regs[31][11] ),
    .S(_02770_),
    .X(_02879_));
 sky130_fd_sc_hd__mux2_1 _08461_ (.A0(\regs[28][11] ),
    .A1(\regs[29][11] ),
    .S(_02395_),
    .X(_02880_));
 sky130_fd_sc_hd__a21o_1 _08462_ (.A1(_02394_),
    .A2(_02880_),
    .B1(_02538_),
    .X(_02881_));
 sky130_fd_sc_hd__a21o_1 _08463_ (.A1(_02299_),
    .A2(_02879_),
    .B1(_02881_),
    .X(_02882_));
 sky130_fd_sc_hd__a31o_1 _08464_ (.A1(_02291_),
    .A2(_02878_),
    .A3(_02882_),
    .B1(_02399_),
    .X(_02883_));
 sky130_fd_sc_hd__a21o_1 _08465_ (.A1(_02366_),
    .A2(_02874_),
    .B1(_02883_),
    .X(_02884_));
 sky130_fd_sc_hd__o221a_1 _08466_ (.A1(_01749_),
    .A2(_02754_),
    .B1(_02709_),
    .B2(_02871_),
    .C1(_02884_),
    .X(_01419_));
 sky130_fd_sc_hd__mux4_1 _08467_ (.A0(\regs[12][10] ),
    .A1(\regs[13][10] ),
    .A2(\regs[14][10] ),
    .A3(\regs[15][10] ),
    .S0(_02340_),
    .S1(_02343_),
    .X(_02885_));
 sky130_fd_sc_hd__or2_1 _08468_ (.A(_02330_),
    .B(_02885_),
    .X(_02886_));
 sky130_fd_sc_hd__mux4_1 _08469_ (.A0(\regs[8][10] ),
    .A1(\regs[9][10] ),
    .A2(\regs[10][10] ),
    .A3(\regs[11][10] ),
    .S0(_02371_),
    .S1(_02402_),
    .X(_02887_));
 sky130_fd_sc_hd__o21a_1 _08470_ (.A1(_02515_),
    .A2(_02887_),
    .B1(_02468_),
    .X(_02888_));
 sky130_fd_sc_hd__mux4_1 _08471_ (.A0(\regs[0][10] ),
    .A1(\regs[1][10] ),
    .A2(\regs[2][10] ),
    .A3(\regs[3][10] ),
    .S0(_02340_),
    .S1(_02336_),
    .X(_02889_));
 sky130_fd_sc_hd__mux4_1 _08472_ (.A0(\regs[4][10] ),
    .A1(\regs[5][10] ),
    .A2(\regs[6][10] ),
    .A3(\regs[7][10] ),
    .S0(_02445_),
    .S1(_02336_),
    .X(_02890_));
 sky130_fd_sc_hd__mux2_1 _08473_ (.A0(_02889_),
    .A1(_02890_),
    .S(_02550_),
    .X(_02891_));
 sky130_fd_sc_hd__a22o_1 _08474_ (.A1(_02886_),
    .A2(_02888_),
    .B1(_02891_),
    .B2(_02362_),
    .X(_02892_));
 sky130_fd_sc_hd__mux4_1 _08475_ (.A0(\regs[16][10] ),
    .A1(\regs[17][10] ),
    .A2(\regs[18][10] ),
    .A3(\regs[19][10] ),
    .S0(_02303_),
    .S1(_02555_),
    .X(_02893_));
 sky130_fd_sc_hd__mux4_1 _08476_ (.A0(\regs[20][10] ),
    .A1(\regs[21][10] ),
    .A2(\regs[22][10] ),
    .A3(\regs[23][10] ),
    .S0(_02303_),
    .S1(_02555_),
    .X(_02894_));
 sky130_fd_sc_hd__mux2_1 _08477_ (.A0(_02893_),
    .A1(_02894_),
    .S(_02294_),
    .X(_02895_));
 sky130_fd_sc_hd__mux2_1 _08478_ (.A0(\regs[30][10] ),
    .A1(\regs[31][10] ),
    .S(_02349_),
    .X(_02896_));
 sky130_fd_sc_hd__mux2_1 _08479_ (.A0(\regs[28][10] ),
    .A1(\regs[29][10] ),
    .S(_02348_),
    .X(_02897_));
 sky130_fd_sc_hd__a21o_1 _08480_ (.A1(_02387_),
    .A2(_02897_),
    .B1(_02418_),
    .X(_02898_));
 sky130_fd_sc_hd__a21o_1 _08481_ (.A1(_02298_),
    .A2(_02896_),
    .B1(_02898_),
    .X(_02899_));
 sky130_fd_sc_hd__or2b_1 _08482_ (.A(\regs[27][10] ),
    .B_N(_02445_),
    .X(_02900_));
 sky130_fd_sc_hd__o21a_1 _08483_ (.A1(_02333_),
    .A2(\regs[26][10] ),
    .B1(_02367_),
    .X(_02901_));
 sky130_fd_sc_hd__mux2_1 _08484_ (.A0(\regs[24][10] ),
    .A1(\regs[25][10] ),
    .S(_02458_),
    .X(_02902_));
 sky130_fd_sc_hd__a221o_1 _08485_ (.A1(_02900_),
    .A2(_02901_),
    .B1(_02902_),
    .B2(_02388_),
    .C1(_02358_),
    .X(_02903_));
 sky130_fd_sc_hd__a31o_1 _08486_ (.A1(_02290_),
    .A2(_02899_),
    .A3(_02903_),
    .B1(_02285_),
    .X(_02904_));
 sky130_fd_sc_hd__a21o_1 _08487_ (.A1(_02365_),
    .A2(_02895_),
    .B1(_02904_),
    .X(_02905_));
 sky130_fd_sc_hd__o211a_1 _08488_ (.A1(_02433_),
    .A2(_02892_),
    .B1(_02905_),
    .C1(_02254_),
    .X(_02906_));
 sky130_fd_sc_hd__a21o_1 _08489_ (.A1(_01877_),
    .A2(_02543_),
    .B1(_02906_),
    .X(_01418_));
 sky130_fd_sc_hd__mux4_1 _08490_ (.A0(\regs[12][9] ),
    .A1(\regs[13][9] ),
    .A2(\regs[14][9] ),
    .A3(\regs[15][9] ),
    .S0(_02350_),
    .S1(_02643_),
    .X(_02907_));
 sky130_fd_sc_hd__or2_1 _08491_ (.A(_02620_),
    .B(_02907_),
    .X(_02908_));
 sky130_fd_sc_hd__mux4_1 _08492_ (.A0(\regs[8][9] ),
    .A1(\regs[9][9] ),
    .A2(\regs[10][9] ),
    .A3(\regs[11][9] ),
    .S0(_02575_),
    .S1(_02576_),
    .X(_02909_));
 sky130_fd_sc_hd__o21a_1 _08493_ (.A1(_02623_),
    .A2(_02909_),
    .B1(_02586_),
    .X(_02910_));
 sky130_fd_sc_hd__mux4_1 _08494_ (.A0(\regs[0][9] ),
    .A1(\regs[1][9] ),
    .A2(\regs[2][9] ),
    .A3(\regs[3][9] ),
    .S0(_02523_),
    .S1(_02356_),
    .X(_02911_));
 sky130_fd_sc_hd__mux4_1 _08495_ (.A0(\regs[4][9] ),
    .A1(\regs[5][9] ),
    .A2(\regs[6][9] ),
    .A3(\regs[7][9] ),
    .S0(_02392_),
    .S1(_02715_),
    .X(_02912_));
 sky130_fd_sc_hd__mux2_1 _08496_ (.A0(_02911_),
    .A1(_02912_),
    .S(_02526_),
    .X(_02913_));
 sky130_fd_sc_hd__a22o_2 _08497_ (.A1(_02908_),
    .A2(_02910_),
    .B1(_02913_),
    .B2(_02569_),
    .X(_02914_));
 sky130_fd_sc_hd__mux4_1 _08498_ (.A0(\regs[20][9] ),
    .A1(\regs[21][9] ),
    .A2(\regs[22][9] ),
    .A3(\regs[23][9] ),
    .S0(_02446_),
    .S1(_02450_),
    .X(_02915_));
 sky130_fd_sc_hd__mux4_1 _08499_ (.A0(\regs[16][9] ),
    .A1(\regs[17][9] ),
    .A2(\regs[18][9] ),
    .A3(\regs[19][9] ),
    .S0(_02449_),
    .S1(_02337_),
    .X(_02916_));
 sky130_fd_sc_hd__mux2_1 _08500_ (.A0(_02915_),
    .A1(_02916_),
    .S(_02452_),
    .X(_02917_));
 sky130_fd_sc_hd__mux2_1 _08501_ (.A0(\regs[30][9] ),
    .A1(\regs[31][9] ),
    .S(_02455_),
    .X(_02918_));
 sky130_fd_sc_hd__and2_1 _08502_ (.A(_02454_),
    .B(_02918_),
    .X(_02919_));
 sky130_fd_sc_hd__mux2_1 _08503_ (.A0(\regs[28][9] ),
    .A1(\regs[29][9] ),
    .S(_02587_),
    .X(_02920_));
 sky130_fd_sc_hd__a21o_1 _08504_ (.A1(_02389_),
    .A2(_02920_),
    .B1(_02422_),
    .X(_02921_));
 sky130_fd_sc_hd__or2b_1 _08505_ (.A(\regs[27][9] ),
    .B_N(_02770_),
    .X(_02922_));
 sky130_fd_sc_hd__o21a_1 _08506_ (.A1(_02770_),
    .A2(\regs[26][9] ),
    .B1(_02368_),
    .X(_02923_));
 sky130_fd_sc_hd__mux2_1 _08507_ (.A0(\regs[24][9] ),
    .A1(\regs[25][9] ),
    .S(_02587_),
    .X(_02924_));
 sky130_fd_sc_hd__a221o_1 _08508_ (.A1(_02922_),
    .A2(_02923_),
    .B1(_02924_),
    .B2(_02466_),
    .C1(_02294_),
    .X(_02925_));
 sky130_fd_sc_hd__o211a_1 _08509_ (.A1(_02919_),
    .A2(_02921_),
    .B1(_02469_),
    .C1(_02925_),
    .X(_02926_));
 sky130_fd_sc_hd__a211o_2 _08510_ (.A1(_02582_),
    .A2(_02917_),
    .B1(_02926_),
    .C1(_02471_),
    .X(_02927_));
 sky130_fd_sc_hd__o221a_1 _08511_ (.A1(_01752_),
    .A2(_02754_),
    .B1(_02709_),
    .B2(_02914_),
    .C1(_02927_),
    .X(_01417_));
 sky130_fd_sc_hd__mux2_1 _08512_ (.A0(\regs[30][8] ),
    .A1(\regs[31][8] ),
    .S(_02403_),
    .X(_02928_));
 sky130_fd_sc_hd__and2_1 _08513_ (.A(_02402_),
    .B(_02928_),
    .X(_02929_));
 sky130_fd_sc_hd__mux2_1 _08514_ (.A0(\regs[28][8] ),
    .A1(\regs[29][8] ),
    .S(_02403_),
    .X(_02930_));
 sky130_fd_sc_hd__a21o_1 _08515_ (.A1(_02413_),
    .A2(_02930_),
    .B1(_02408_),
    .X(_02931_));
 sky130_fd_sc_hd__or2b_1 _08516_ (.A(\regs[27][8] ),
    .B_N(_02380_),
    .X(_02932_));
 sky130_fd_sc_hd__o21a_1 _08517_ (.A1(_02406_),
    .A2(\regs[26][8] ),
    .B1(_02335_),
    .X(_02933_));
 sky130_fd_sc_hd__mux2_1 _08518_ (.A0(\regs[24][8] ),
    .A1(\regs[25][8] ),
    .S(_02302_),
    .X(_02934_));
 sky130_fd_sc_hd__a221o_1 _08519_ (.A1(_02932_),
    .A2(_02933_),
    .B1(_02934_),
    .B2(_02387_),
    .C1(net10),
    .X(_02935_));
 sky130_fd_sc_hd__o211a_1 _08520_ (.A1(_02929_),
    .A2(_02931_),
    .B1(_02935_),
    .C1(_02289_),
    .X(_02936_));
 sky130_fd_sc_hd__mux4_1 _08521_ (.A0(\regs[16][8] ),
    .A1(\regs[17][8] ),
    .A2(\regs[18][8] ),
    .A3(\regs[19][8] ),
    .S0(_02349_),
    .S1(_02351_),
    .X(_02937_));
 sky130_fd_sc_hd__mux4_1 _08522_ (.A0(\regs[20][8] ),
    .A1(\regs[21][8] ),
    .A2(\regs[22][8] ),
    .A3(\regs[23][8] ),
    .S0(_02301_),
    .S1(_02335_),
    .X(_02938_));
 sky130_fd_sc_hd__or2_1 _08523_ (.A(_02418_),
    .B(_02938_),
    .X(_02939_));
 sky130_fd_sc_hd__o211a_1 _08524_ (.A1(_02375_),
    .A2(_02937_),
    .B1(_02939_),
    .C1(_02361_),
    .X(_02940_));
 sky130_fd_sc_hd__mux4_1 _08525_ (.A0(\regs[12][8] ),
    .A1(\regs[13][8] ),
    .A2(\regs[14][8] ),
    .A3(\regs[15][8] ),
    .S0(_02371_),
    .S1(_02423_),
    .X(_02941_));
 sky130_fd_sc_hd__mux4_1 _08526_ (.A0(\regs[8][8] ),
    .A1(\regs[9][8] ),
    .A2(\regs[10][8] ),
    .A3(\regs[11][8] ),
    .S0(_02428_),
    .S1(_02429_),
    .X(_02942_));
 sky130_fd_sc_hd__or2_1 _08527_ (.A(_02293_),
    .B(_02942_),
    .X(_02943_));
 sky130_fd_sc_hd__o211a_1 _08528_ (.A1(_02422_),
    .A2(_02941_),
    .B1(_02943_),
    .C1(_02468_),
    .X(_02944_));
 sky130_fd_sc_hd__mux4_1 _08529_ (.A0(\regs[0][8] ),
    .A1(\regs[1][8] ),
    .A2(\regs[2][8] ),
    .A3(\regs[3][8] ),
    .S0(_02428_),
    .S1(_02429_),
    .X(_02945_));
 sky130_fd_sc_hd__mux4_1 _08530_ (.A0(\regs[4][8] ),
    .A1(\regs[5][8] ),
    .A2(\regs[6][8] ),
    .A3(\regs[7][8] ),
    .S0(_02332_),
    .S1(_02342_),
    .X(_02946_));
 sky130_fd_sc_hd__mux2_1 _08531_ (.A0(_02945_),
    .A1(_02946_),
    .S(_02414_),
    .X(_02947_));
 sky130_fd_sc_hd__a21o_1 _08532_ (.A1(_02361_),
    .A2(_02947_),
    .B1(net12),
    .X(_02948_));
 sky130_fd_sc_hd__o32a_2 _08533_ (.A1(_02286_),
    .A2(_02936_),
    .A3(_02940_),
    .B1(_02944_),
    .B2(_02948_),
    .X(_02949_));
 sky130_fd_sc_hd__mux2_1 _08534_ (.A0(\leorv32_alu.input1[8] ),
    .A1(_02949_),
    .S(_02324_),
    .X(_02950_));
 sky130_fd_sc_hd__clkbuf_1 _08535_ (.A(_02950_),
    .X(_01416_));
 sky130_fd_sc_hd__mux4_1 _08536_ (.A0(\regs[0][7] ),
    .A1(\regs[1][7] ),
    .A2(\regs[2][7] ),
    .A3(\regs[3][7] ),
    .S0(_02462_),
    .S1(_02298_),
    .X(_02951_));
 sky130_fd_sc_hd__mux4_1 _08537_ (.A0(\regs[4][7] ),
    .A1(\regs[5][7] ),
    .A2(\regs[6][7] ),
    .A3(\regs[7][7] ),
    .S0(_02571_),
    .S1(_02572_),
    .X(_02952_));
 sky130_fd_sc_hd__mux2_1 _08538_ (.A0(_02951_),
    .A1(_02952_),
    .S(_02390_),
    .X(_02953_));
 sky130_fd_sc_hd__mux4_1 _08539_ (.A0(\regs[8][7] ),
    .A1(\regs[9][7] ),
    .A2(\regs[10][7] ),
    .A3(\regs[11][7] ),
    .S0(_02446_),
    .S1(_02447_),
    .X(_02954_));
 sky130_fd_sc_hd__or2_1 _08540_ (.A(_02623_),
    .B(_02954_),
    .X(_02955_));
 sky130_fd_sc_hd__mux4_1 _08541_ (.A0(\regs[12][7] ),
    .A1(\regs[13][7] ),
    .A2(\regs[14][7] ),
    .A3(\regs[15][7] ),
    .S0(_02341_),
    .S1(_02344_),
    .X(_02956_));
 sky130_fd_sc_hd__o21a_1 _08542_ (.A1(_02331_),
    .A2(_02956_),
    .B1(_02469_),
    .X(_02957_));
 sky130_fd_sc_hd__a22o_2 _08543_ (.A1(_02569_),
    .A2(_02953_),
    .B1(_02955_),
    .B2(_02957_),
    .X(_02958_));
 sky130_fd_sc_hd__mux4_1 _08544_ (.A0(\regs[16][7] ),
    .A1(\regs[17][7] ),
    .A2(\regs[18][7] ),
    .A3(\regs[19][7] ),
    .S0(_02449_),
    .S1(_02450_),
    .X(_02959_));
 sky130_fd_sc_hd__mux4_1 _08545_ (.A0(\regs[20][7] ),
    .A1(\regs[21][7] ),
    .A2(\regs[22][7] ),
    .A3(\regs[23][7] ),
    .S0(_02378_),
    .S1(_02337_),
    .X(_02960_));
 sky130_fd_sc_hd__mux2_1 _08546_ (.A0(_02959_),
    .A1(_02960_),
    .S(_02359_),
    .X(_02961_));
 sky130_fd_sc_hd__mux2_1 _08547_ (.A0(\regs[30][7] ),
    .A1(\regs[31][7] ),
    .S(_02587_),
    .X(_02962_));
 sky130_fd_sc_hd__mux2_1 _08548_ (.A0(\regs[28][7] ),
    .A1(\regs[29][7] ),
    .S(_02354_),
    .X(_02963_));
 sky130_fd_sc_hd__a21o_1 _08549_ (.A1(_02394_),
    .A2(_02963_),
    .B1(_02538_),
    .X(_02964_));
 sky130_fd_sc_hd__a21o_1 _08550_ (.A1(_02454_),
    .A2(_02962_),
    .B1(_02964_),
    .X(_02965_));
 sky130_fd_sc_hd__or2b_1 _08551_ (.A(\regs[27][7] ),
    .B_N(_02592_),
    .X(_02966_));
 sky130_fd_sc_hd__o21a_1 _08552_ (.A1(_02384_),
    .A2(\regs[26][7] ),
    .B1(_02423_),
    .X(_02967_));
 sky130_fd_sc_hd__mux2_1 _08553_ (.A0(\regs[24][7] ),
    .A1(\regs[25][7] ),
    .S(_02553_),
    .X(_02968_));
 sky130_fd_sc_hd__a221o_1 _08554_ (.A1(_02966_),
    .A2(_02967_),
    .B1(_02968_),
    .B2(_02508_),
    .C1(_02550_),
    .X(_02969_));
 sky130_fd_sc_hd__and3_1 _08555_ (.A(_02586_),
    .B(_02965_),
    .C(_02969_),
    .X(_02970_));
 sky130_fd_sc_hd__a211o_1 _08556_ (.A1(_02582_),
    .A2(_02961_),
    .B1(_02970_),
    .C1(_02471_),
    .X(_02971_));
 sky130_fd_sc_hd__o221a_1 _08557_ (.A1(_01784_),
    .A2(_02754_),
    .B1(_02709_),
    .B2(_02958_),
    .C1(_02971_),
    .X(_01415_));
 sky130_fd_sc_hd__mux4_1 _08558_ (.A0(\regs[16][6] ),
    .A1(\regs[17][6] ),
    .A2(\regs[18][6] ),
    .A3(\regs[19][6] ),
    .S0(_02770_),
    .S1(_02715_),
    .X(_02972_));
 sky130_fd_sc_hd__mux4_1 _08559_ (.A0(\regs[20][6] ),
    .A1(\regs[21][6] ),
    .A2(\regs[22][6] ),
    .A3(\regs[23][6] ),
    .S0(_02770_),
    .S1(_02715_),
    .X(_02973_));
 sky130_fd_sc_hd__mux2_1 _08560_ (.A0(_02972_),
    .A1(_02973_),
    .S(_02390_),
    .X(_02974_));
 sky130_fd_sc_hd__mux2_1 _08561_ (.A0(\regs[30][6] ),
    .A1(\regs[31][6] ),
    .S(_02455_),
    .X(_02975_));
 sky130_fd_sc_hd__and2_1 _08562_ (.A(_02369_),
    .B(_02975_),
    .X(_02976_));
 sky130_fd_sc_hd__mux2_1 _08563_ (.A0(\regs[28][6] ),
    .A1(\regs[29][6] ),
    .S(_02455_),
    .X(_02977_));
 sky130_fd_sc_hd__a21o_1 _08564_ (.A1(_02466_),
    .A2(_02977_),
    .B1(_02422_),
    .X(_02978_));
 sky130_fd_sc_hd__or2b_1 _08565_ (.A(\regs[27][6] ),
    .B_N(_02592_),
    .X(_02979_));
 sky130_fd_sc_hd__o21a_1 _08566_ (.A1(_02592_),
    .A2(\regs[26][6] ),
    .B1(_02555_),
    .X(_02980_));
 sky130_fd_sc_hd__mux2_1 _08567_ (.A0(\regs[24][6] ),
    .A1(\regs[25][6] ),
    .S(_02553_),
    .X(_02981_));
 sky130_fd_sc_hd__a221o_1 _08568_ (.A1(_02979_),
    .A2(_02980_),
    .B1(_02981_),
    .B2(_02508_),
    .C1(_02550_),
    .X(_02982_));
 sky130_fd_sc_hd__o211a_1 _08569_ (.A1(_02976_),
    .A2(_02978_),
    .B1(_02982_),
    .C1(_02346_),
    .X(_02983_));
 sky130_fd_sc_hd__a211o_1 _08570_ (.A1(_02363_),
    .A2(_02974_),
    .B1(_02983_),
    .C1(_02286_),
    .X(_02984_));
 sky130_fd_sc_hd__mux4_1 _08571_ (.A0(\regs[12][6] ),
    .A1(\regs[13][6] ),
    .A2(\regs[14][6] ),
    .A3(\regs[15][6] ),
    .S0(_02462_),
    .S1(_02298_),
    .X(_02985_));
 sky130_fd_sc_hd__or2_1 _08572_ (.A(_02452_),
    .B(_02985_),
    .X(_02986_));
 sky130_fd_sc_hd__mux4_1 _08573_ (.A0(\regs[8][6] ),
    .A1(\regs[9][6] ),
    .A2(\regs[10][6] ),
    .A3(\regs[11][6] ),
    .S0(_02350_),
    .S1(_02643_),
    .X(_02987_));
 sky130_fd_sc_hd__o21a_1 _08574_ (.A1(_02359_),
    .A2(_02987_),
    .B1(_02290_),
    .X(_02988_));
 sky130_fd_sc_hd__mux4_1 _08575_ (.A0(\regs[0][6] ),
    .A1(\regs[1][6] ),
    .A2(\regs[2][6] ),
    .A3(\regs[3][6] ),
    .S0(_02571_),
    .S1(_02382_),
    .X(_02989_));
 sky130_fd_sc_hd__mux4_1 _08576_ (.A0(\regs[4][6] ),
    .A1(\regs[5][6] ),
    .A2(\regs[6][6] ),
    .A3(\regs[7][6] ),
    .S0(_02592_),
    .S1(_02382_),
    .X(_02990_));
 sky130_fd_sc_hd__mux2_1 _08577_ (.A0(_02989_),
    .A1(_02990_),
    .S(_02390_),
    .X(_02991_));
 sky130_fd_sc_hd__a221o_2 _08578_ (.A1(_02986_),
    .A2(_02988_),
    .B1(_02991_),
    .B2(_02365_),
    .C1(_02433_),
    .X(_02992_));
 sky130_fd_sc_hd__buf_4 _08579_ (.A(_02253_),
    .X(_02993_));
 sky130_fd_sc_hd__nor2_1 _08580_ (.A(_01767_),
    .B(_02993_),
    .Y(_02994_));
 sky130_fd_sc_hd__a31o_1 _08581_ (.A1(_00001_),
    .A2(_02984_),
    .A3(_02992_),
    .B1(_02994_),
    .X(_01414_));
 sky130_fd_sc_hd__mux2_1 _08582_ (.A0(\regs[30][5] ),
    .A1(\regs[31][5] ),
    .S(_02403_),
    .X(_02995_));
 sky130_fd_sc_hd__and2_1 _08583_ (.A(_02402_),
    .B(_02995_),
    .X(_02996_));
 sky130_fd_sc_hd__mux2_1 _08584_ (.A0(\regs[28][5] ),
    .A1(\regs[29][5] ),
    .S(_02403_),
    .X(_02997_));
 sky130_fd_sc_hd__a21o_1 _08585_ (.A1(_02413_),
    .A2(_02997_),
    .B1(_02408_),
    .X(_02998_));
 sky130_fd_sc_hd__or2b_1 _08586_ (.A(\regs[27][5] ),
    .B_N(_02380_),
    .X(_02999_));
 sky130_fd_sc_hd__o21a_1 _08587_ (.A1(_02406_),
    .A2(\regs[26][5] ),
    .B1(_02335_),
    .X(_03000_));
 sky130_fd_sc_hd__mux2_1 _08588_ (.A0(\regs[24][5] ),
    .A1(\regs[25][5] ),
    .S(_02302_),
    .X(_03001_));
 sky130_fd_sc_hd__a221o_1 _08589_ (.A1(_02999_),
    .A2(_03000_),
    .B1(_03001_),
    .B2(_02387_),
    .C1(net10),
    .X(_03002_));
 sky130_fd_sc_hd__o211a_1 _08590_ (.A1(_02996_),
    .A2(_02998_),
    .B1(_03002_),
    .C1(_02289_),
    .X(_03003_));
 sky130_fd_sc_hd__mux4_1 _08591_ (.A0(\regs[16][5] ),
    .A1(\regs[17][5] ),
    .A2(\regs[18][5] ),
    .A3(\regs[19][5] ),
    .S0(_02349_),
    .S1(_02351_),
    .X(_03004_));
 sky130_fd_sc_hd__mux4_1 _08592_ (.A0(\regs[20][5] ),
    .A1(\regs[21][5] ),
    .A2(\regs[22][5] ),
    .A3(\regs[23][5] ),
    .S0(_02301_),
    .S1(_02335_),
    .X(_03005_));
 sky130_fd_sc_hd__or2_1 _08593_ (.A(_02418_),
    .B(_03005_),
    .X(_03006_));
 sky130_fd_sc_hd__o211a_1 _08594_ (.A1(_02375_),
    .A2(_03004_),
    .B1(_03006_),
    .C1(_02361_),
    .X(_03007_));
 sky130_fd_sc_hd__mux4_1 _08595_ (.A0(\regs[12][5] ),
    .A1(\regs[13][5] ),
    .A2(\regs[14][5] ),
    .A3(\regs[15][5] ),
    .S0(_02371_),
    .S1(_02423_),
    .X(_03008_));
 sky130_fd_sc_hd__mux4_1 _08596_ (.A0(\regs[8][5] ),
    .A1(\regs[9][5] ),
    .A2(\regs[10][5] ),
    .A3(\regs[11][5] ),
    .S0(_02428_),
    .S1(_02429_),
    .X(_03009_));
 sky130_fd_sc_hd__or2_1 _08597_ (.A(_02293_),
    .B(_03009_),
    .X(_03010_));
 sky130_fd_sc_hd__o211a_1 _08598_ (.A1(_02422_),
    .A2(_03008_),
    .B1(_03010_),
    .C1(_02468_),
    .X(_03011_));
 sky130_fd_sc_hd__mux4_1 _08599_ (.A0(\regs[0][5] ),
    .A1(\regs[1][5] ),
    .A2(\regs[2][5] ),
    .A3(\regs[3][5] ),
    .S0(_02332_),
    .S1(_02429_),
    .X(_03012_));
 sky130_fd_sc_hd__mux4_1 _08600_ (.A0(\regs[4][5] ),
    .A1(\regs[5][5] ),
    .A2(\regs[6][5] ),
    .A3(\regs[7][5] ),
    .S0(_02332_),
    .S1(_02342_),
    .X(_03013_));
 sky130_fd_sc_hd__mux2_1 _08601_ (.A0(_03012_),
    .A1(_03013_),
    .S(_02414_),
    .X(_03014_));
 sky130_fd_sc_hd__a21o_1 _08602_ (.A1(_02361_),
    .A2(_03014_),
    .B1(net12),
    .X(_03015_));
 sky130_fd_sc_hd__o32a_2 _08603_ (.A1(_02286_),
    .A2(_03003_),
    .A3(_03007_),
    .B1(_03011_),
    .B2(_03015_),
    .X(_03016_));
 sky130_fd_sc_hd__mux2_1 _08604_ (.A0(\leorv32_alu.input1[5] ),
    .A1(_03016_),
    .S(_02324_),
    .X(_03017_));
 sky130_fd_sc_hd__clkbuf_1 _08605_ (.A(_03017_),
    .X(_01413_));
 sky130_fd_sc_hd__mux4_1 _08606_ (.A0(\regs[12][4] ),
    .A1(\regs[13][4] ),
    .A2(\regs[14][4] ),
    .A3(\regs[15][4] ),
    .S0(_02340_),
    .S1(_02343_),
    .X(_03018_));
 sky130_fd_sc_hd__or2_1 _08607_ (.A(_02330_),
    .B(_03018_),
    .X(_03019_));
 sky130_fd_sc_hd__mux4_1 _08608_ (.A0(\regs[8][4] ),
    .A1(\regs[9][4] ),
    .A2(\regs[10][4] ),
    .A3(\regs[11][4] ),
    .S0(_02371_),
    .S1(_02402_),
    .X(_03020_));
 sky130_fd_sc_hd__o21a_1 _08609_ (.A1(_02294_),
    .A2(_03020_),
    .B1(_02468_),
    .X(_03021_));
 sky130_fd_sc_hd__mux4_1 _08610_ (.A0(\regs[0][4] ),
    .A1(\regs[1][4] ),
    .A2(\regs[2][4] ),
    .A3(\regs[3][4] ),
    .S0(_02340_),
    .S1(_02336_),
    .X(_03022_));
 sky130_fd_sc_hd__mux4_1 _08611_ (.A0(\regs[4][4] ),
    .A1(\regs[5][4] ),
    .A2(\regs[6][4] ),
    .A3(\regs[7][4] ),
    .S0(_02445_),
    .S1(_02336_),
    .X(_03023_));
 sky130_fd_sc_hd__mux2_1 _08612_ (.A0(_03022_),
    .A1(_03023_),
    .S(_02358_),
    .X(_03024_));
 sky130_fd_sc_hd__a22o_1 _08613_ (.A1(_03019_),
    .A2(_03021_),
    .B1(_03024_),
    .B2(_02362_),
    .X(_03025_));
 sky130_fd_sc_hd__mux4_1 _08614_ (.A0(\regs[16][4] ),
    .A1(\regs[17][4] ),
    .A2(\regs[18][4] ),
    .A3(\regs[19][4] ),
    .S0(_02303_),
    .S1(_02555_),
    .X(_03026_));
 sky130_fd_sc_hd__mux4_1 _08615_ (.A0(\regs[20][4] ),
    .A1(\regs[21][4] ),
    .A2(\regs[22][4] ),
    .A3(\regs[23][4] ),
    .S0(_02303_),
    .S1(_02555_),
    .X(_03027_));
 sky130_fd_sc_hd__mux2_1 _08616_ (.A0(_03026_),
    .A1(_03027_),
    .S(_02375_),
    .X(_03028_));
 sky130_fd_sc_hd__mux2_1 _08617_ (.A0(\regs[30][4] ),
    .A1(\regs[31][4] ),
    .S(_02349_),
    .X(_03029_));
 sky130_fd_sc_hd__mux2_1 _08618_ (.A0(\regs[28][4] ),
    .A1(\regs[29][4] ),
    .S(_02348_),
    .X(_03030_));
 sky130_fd_sc_hd__a21o_1 _08619_ (.A1(_02387_),
    .A2(_03030_),
    .B1(_02418_),
    .X(_03031_));
 sky130_fd_sc_hd__a21o_1 _08620_ (.A1(_02298_),
    .A2(_03029_),
    .B1(_03031_),
    .X(_03032_));
 sky130_fd_sc_hd__or2b_1 _08621_ (.A(\regs[27][4] ),
    .B_N(_02445_),
    .X(_03033_));
 sky130_fd_sc_hd__o21a_1 _08622_ (.A1(_02333_),
    .A2(\regs[26][4] ),
    .B1(_02367_),
    .X(_03034_));
 sky130_fd_sc_hd__mux2_1 _08623_ (.A0(\regs[24][4] ),
    .A1(\regs[25][4] ),
    .S(_02458_),
    .X(_03035_));
 sky130_fd_sc_hd__a221o_1 _08624_ (.A1(_03033_),
    .A2(_03034_),
    .B1(_03035_),
    .B2(_02388_),
    .C1(_02358_),
    .X(_03036_));
 sky130_fd_sc_hd__a31o_1 _08625_ (.A1(_02290_),
    .A2(_03032_),
    .A3(_03036_),
    .B1(_02285_),
    .X(_03037_));
 sky130_fd_sc_hd__a21o_1 _08626_ (.A1(_02365_),
    .A2(_03028_),
    .B1(_03037_),
    .X(_03038_));
 sky130_fd_sc_hd__o211a_2 _08627_ (.A1(_02433_),
    .A2(_03025_),
    .B1(_03038_),
    .C1(_02254_),
    .X(_03039_));
 sky130_fd_sc_hd__a21o_1 _08628_ (.A1(_01764_),
    .A2(_02543_),
    .B1(_03039_),
    .X(_01412_));
 sky130_fd_sc_hd__mux4_1 _08629_ (.A0(\regs[4][3] ),
    .A1(\regs[5][3] ),
    .A2(\regs[6][3] ),
    .A3(\regs[7][3] ),
    .S0(_02462_),
    .S1(_02572_),
    .X(_03040_));
 sky130_fd_sc_hd__mux4_1 _08630_ (.A0(\regs[0][3] ),
    .A1(\regs[1][3] ),
    .A2(\regs[2][3] ),
    .A3(\regs[3][3] ),
    .S0(_02571_),
    .S1(_02572_),
    .X(_03041_));
 sky130_fd_sc_hd__mux2_1 _08631_ (.A0(_03040_),
    .A1(_03041_),
    .S(_02452_),
    .X(_03042_));
 sky130_fd_sc_hd__mux4_1 _08632_ (.A0(\regs[12][3] ),
    .A1(\regs[13][3] ),
    .A2(\regs[14][3] ),
    .A3(\regs[15][3] ),
    .S0(_02446_),
    .S1(_02447_),
    .X(_03043_));
 sky130_fd_sc_hd__or2_1 _08633_ (.A(_02331_),
    .B(_03043_),
    .X(_03044_));
 sky130_fd_sc_hd__mux4_1 _08634_ (.A0(\regs[8][3] ),
    .A1(\regs[9][3] ),
    .A2(\regs[10][3] ),
    .A3(\regs[11][3] ),
    .S0(_02341_),
    .S1(_02344_),
    .X(_03045_));
 sky130_fd_sc_hd__o21a_1 _08635_ (.A1(_02295_),
    .A2(_03045_),
    .B1(_02469_),
    .X(_03046_));
 sky130_fd_sc_hd__a22o_2 _08636_ (.A1(_02569_),
    .A2(_03042_),
    .B1(_03044_),
    .B2(_03046_),
    .X(_03047_));
 sky130_fd_sc_hd__mux4_1 _08637_ (.A0(\regs[16][3] ),
    .A1(\regs[17][3] ),
    .A2(\regs[18][3] ),
    .A3(\regs[19][3] ),
    .S0(_02449_),
    .S1(_02450_),
    .X(_03048_));
 sky130_fd_sc_hd__mux4_1 _08638_ (.A0(\regs[20][3] ),
    .A1(\regs[21][3] ),
    .A2(\regs[22][3] ),
    .A3(\regs[23][3] ),
    .S0(_02378_),
    .S1(_02337_),
    .X(_03049_));
 sky130_fd_sc_hd__mux2_1 _08639_ (.A0(_03048_),
    .A1(_03049_),
    .S(_02359_),
    .X(_03050_));
 sky130_fd_sc_hd__mux2_1 _08640_ (.A0(\regs[30][3] ),
    .A1(\regs[31][3] ),
    .S(_02587_),
    .X(_03051_));
 sky130_fd_sc_hd__mux2_1 _08641_ (.A0(\regs[28][3] ),
    .A1(\regs[29][3] ),
    .S(_02458_),
    .X(_03052_));
 sky130_fd_sc_hd__a21o_1 _08642_ (.A1(_02388_),
    .A2(_03052_),
    .B1(_02538_),
    .X(_03053_));
 sky130_fd_sc_hd__a21o_1 _08643_ (.A1(_02454_),
    .A2(_03051_),
    .B1(_03053_),
    .X(_03054_));
 sky130_fd_sc_hd__or2b_1 _08644_ (.A(\regs[27][3] ),
    .B_N(_02592_),
    .X(_03055_));
 sky130_fd_sc_hd__o21a_1 _08645_ (.A1(_02384_),
    .A2(\regs[26][3] ),
    .B1(_02423_),
    .X(_03056_));
 sky130_fd_sc_hd__mux2_1 _08646_ (.A0(\regs[24][3] ),
    .A1(\regs[25][3] ),
    .S(_02553_),
    .X(_03057_));
 sky130_fd_sc_hd__a221o_1 _08647_ (.A1(_03055_),
    .A2(_03056_),
    .B1(_03057_),
    .B2(_02508_),
    .C1(_02550_),
    .X(_03058_));
 sky130_fd_sc_hd__and3_1 _08648_ (.A(_02586_),
    .B(_03054_),
    .C(_03058_),
    .X(_03059_));
 sky130_fd_sc_hd__a211o_2 _08649_ (.A1(_02582_),
    .A2(_03050_),
    .B1(_03059_),
    .C1(_02471_),
    .X(_03060_));
 sky130_fd_sc_hd__o221a_1 _08650_ (.A1(_01898_),
    .A2(_02754_),
    .B1(_02709_),
    .B2(_03047_),
    .C1(_03060_),
    .X(_01411_));
 sky130_fd_sc_hd__mux4_1 _08651_ (.A0(\regs[0][2] ),
    .A1(\regs[1][2] ),
    .A2(\regs[2][2] ),
    .A3(\regs[3][2] ),
    .S0(_02571_),
    .S1(_02572_),
    .X(_03061_));
 sky130_fd_sc_hd__mux4_1 _08652_ (.A0(\regs[4][2] ),
    .A1(\regs[5][2] ),
    .A2(\regs[6][2] ),
    .A3(\regs[7][2] ),
    .S0(_02571_),
    .S1(_02572_),
    .X(_03062_));
 sky130_fd_sc_hd__mux2_1 _08653_ (.A0(_03061_),
    .A1(_03062_),
    .S(_02390_),
    .X(_03063_));
 sky130_fd_sc_hd__mux4_1 _08654_ (.A0(\regs[12][2] ),
    .A1(\regs[13][2] ),
    .A2(\regs[14][2] ),
    .A3(\regs[15][2] ),
    .S0(_02446_),
    .S1(_02447_),
    .X(_03064_));
 sky130_fd_sc_hd__or2_1 _08655_ (.A(_02331_),
    .B(_03064_),
    .X(_03065_));
 sky130_fd_sc_hd__mux4_1 _08656_ (.A0(\regs[8][2] ),
    .A1(\regs[9][2] ),
    .A2(\regs[10][2] ),
    .A3(\regs[11][2] ),
    .S0(_02341_),
    .S1(_02344_),
    .X(_03066_));
 sky130_fd_sc_hd__o21a_1 _08657_ (.A1(_02295_),
    .A2(_03066_),
    .B1(_02469_),
    .X(_03067_));
 sky130_fd_sc_hd__a22o_2 _08658_ (.A1(_02569_),
    .A2(_03063_),
    .B1(_03065_),
    .B2(_03067_),
    .X(_03068_));
 sky130_fd_sc_hd__mux4_1 _08659_ (.A0(\regs[16][2] ),
    .A1(\regs[17][2] ),
    .A2(\regs[18][2] ),
    .A3(\regs[19][2] ),
    .S0(_02449_),
    .S1(_02450_),
    .X(_03069_));
 sky130_fd_sc_hd__mux4_1 _08660_ (.A0(\regs[20][2] ),
    .A1(\regs[21][2] ),
    .A2(\regs[22][2] ),
    .A3(\regs[23][2] ),
    .S0(_02378_),
    .S1(_02337_),
    .X(_03070_));
 sky130_fd_sc_hd__mux2_1 _08661_ (.A0(_03069_),
    .A1(_03070_),
    .S(_02359_),
    .X(_03071_));
 sky130_fd_sc_hd__mux2_1 _08662_ (.A0(\regs[30][2] ),
    .A1(\regs[31][2] ),
    .S(_02587_),
    .X(_03072_));
 sky130_fd_sc_hd__mux2_1 _08663_ (.A0(\regs[28][2] ),
    .A1(\regs[29][2] ),
    .S(_02458_),
    .X(_03073_));
 sky130_fd_sc_hd__a21o_1 _08664_ (.A1(_02388_),
    .A2(_03073_),
    .B1(_02408_),
    .X(_03074_));
 sky130_fd_sc_hd__a21o_1 _08665_ (.A1(_02454_),
    .A2(_03072_),
    .B1(_03074_),
    .X(_03075_));
 sky130_fd_sc_hd__or2b_1 _08666_ (.A(\regs[27][2] ),
    .B_N(_02384_),
    .X(_03076_));
 sky130_fd_sc_hd__o21a_1 _08667_ (.A1(_02384_),
    .A2(\regs[26][2] ),
    .B1(_02423_),
    .X(_03077_));
 sky130_fd_sc_hd__mux2_1 _08668_ (.A0(\regs[24][2] ),
    .A1(\regs[25][2] ),
    .S(_02553_),
    .X(_03078_));
 sky130_fd_sc_hd__a221o_1 _08669_ (.A1(_03076_),
    .A2(_03077_),
    .B1(_03078_),
    .B2(_02508_),
    .C1(_02550_),
    .X(_03079_));
 sky130_fd_sc_hd__and3_1 _08670_ (.A(_02586_),
    .B(_03075_),
    .C(_03079_),
    .X(_03080_));
 sky130_fd_sc_hd__a211o_2 _08671_ (.A1(_02582_),
    .A2(_03071_),
    .B1(_03080_),
    .C1(_02471_),
    .X(_03081_));
 sky130_fd_sc_hd__o221a_1 _08672_ (.A1(_01901_),
    .A2(_02754_),
    .B1(_02709_),
    .B2(_03068_),
    .C1(_03081_),
    .X(_01410_));
 sky130_fd_sc_hd__mux4_1 _08673_ (.A0(\regs[0][1] ),
    .A1(\regs[1][1] ),
    .A2(\regs[2][1] ),
    .A3(\regs[3][1] ),
    .S0(_02571_),
    .S1(_02572_),
    .X(_03082_));
 sky130_fd_sc_hd__mux4_1 _08674_ (.A0(\regs[4][1] ),
    .A1(\regs[5][1] ),
    .A2(\regs[6][1] ),
    .A3(\regs[7][1] ),
    .S0(_02571_),
    .S1(_02572_),
    .X(_03083_));
 sky130_fd_sc_hd__mux2_1 _08675_ (.A0(_03082_),
    .A1(_03083_),
    .S(_02390_),
    .X(_03084_));
 sky130_fd_sc_hd__mux4_1 _08676_ (.A0(\regs[12][1] ),
    .A1(\regs[13][1] ),
    .A2(\regs[14][1] ),
    .A3(\regs[15][1] ),
    .S0(_02446_),
    .S1(_02447_),
    .X(_03085_));
 sky130_fd_sc_hd__or2_1 _08677_ (.A(_02331_),
    .B(_03085_),
    .X(_03086_));
 sky130_fd_sc_hd__mux4_1 _08678_ (.A0(\regs[8][1] ),
    .A1(\regs[9][1] ),
    .A2(\regs[10][1] ),
    .A3(\regs[11][1] ),
    .S0(_02341_),
    .S1(_02344_),
    .X(_03087_));
 sky130_fd_sc_hd__o21a_1 _08679_ (.A1(_02295_),
    .A2(_03087_),
    .B1(_02469_),
    .X(_03088_));
 sky130_fd_sc_hd__a22o_2 _08680_ (.A1(_02569_),
    .A2(_03084_),
    .B1(_03086_),
    .B2(_03088_),
    .X(_03089_));
 sky130_fd_sc_hd__mux4_1 _08681_ (.A0(\regs[16][1] ),
    .A1(\regs[17][1] ),
    .A2(\regs[18][1] ),
    .A3(\regs[19][1] ),
    .S0(_02449_),
    .S1(_02450_),
    .X(_03090_));
 sky130_fd_sc_hd__mux4_1 _08682_ (.A0(\regs[20][1] ),
    .A1(\regs[21][1] ),
    .A2(\regs[22][1] ),
    .A3(\regs[23][1] ),
    .S0(_02378_),
    .S1(_02337_),
    .X(_03091_));
 sky130_fd_sc_hd__mux2_1 _08683_ (.A0(_03090_),
    .A1(_03091_),
    .S(_02359_),
    .X(_03092_));
 sky130_fd_sc_hd__mux2_1 _08684_ (.A0(\regs[30][1] ),
    .A1(\regs[31][1] ),
    .S(_02587_),
    .X(_03093_));
 sky130_fd_sc_hd__mux2_1 _08685_ (.A0(\regs[28][1] ),
    .A1(\regs[29][1] ),
    .S(_02458_),
    .X(_03094_));
 sky130_fd_sc_hd__a21o_1 _08686_ (.A1(_02388_),
    .A2(_03094_),
    .B1(_02408_),
    .X(_03095_));
 sky130_fd_sc_hd__a21o_1 _08687_ (.A1(_02454_),
    .A2(_03093_),
    .B1(_03095_),
    .X(_03096_));
 sky130_fd_sc_hd__or2b_1 _08688_ (.A(\regs[27][1] ),
    .B_N(_02384_),
    .X(_03097_));
 sky130_fd_sc_hd__o21a_1 _08689_ (.A1(_02384_),
    .A2(\regs[26][1] ),
    .B1(_02423_),
    .X(_03098_));
 sky130_fd_sc_hd__mux2_1 _08690_ (.A0(\regs[24][1] ),
    .A1(\regs[25][1] ),
    .S(_02553_),
    .X(_03099_));
 sky130_fd_sc_hd__a221o_1 _08691_ (.A1(_03097_),
    .A2(_03098_),
    .B1(_03099_),
    .B2(_02508_),
    .C1(_02550_),
    .X(_03100_));
 sky130_fd_sc_hd__and3_1 _08692_ (.A(_02290_),
    .B(_03096_),
    .C(_03100_),
    .X(_03101_));
 sky130_fd_sc_hd__a211o_2 _08693_ (.A1(_02582_),
    .A2(_03092_),
    .B1(_03101_),
    .C1(_02471_),
    .X(_03102_));
 sky130_fd_sc_hd__o221a_1 _08694_ (.A1(_01778_),
    .A2(_02754_),
    .B1(_02709_),
    .B2(_03089_),
    .C1(_03102_),
    .X(_01409_));
 sky130_fd_sc_hd__mux4_1 _08695_ (.A0(\regs[16][0] ),
    .A1(\regs[17][0] ),
    .A2(\regs[18][0] ),
    .A3(\regs[19][0] ),
    .S0(_02371_),
    .S1(_02343_),
    .X(_03103_));
 sky130_fd_sc_hd__mux4_1 _08696_ (.A0(\regs[20][0] ),
    .A1(\regs[21][0] ),
    .A2(\regs[22][0] ),
    .A3(\regs[23][0] ),
    .S0(_02371_),
    .S1(_02343_),
    .X(_03104_));
 sky130_fd_sc_hd__mux2_1 _08697_ (.A0(_03103_),
    .A1(_03104_),
    .S(_02375_),
    .X(_03105_));
 sky130_fd_sc_hd__mux2_1 _08698_ (.A0(\regs[28][0] ),
    .A1(\regs[29][0] ),
    .S(_02354_),
    .X(_03106_));
 sky130_fd_sc_hd__mux2_1 _08699_ (.A0(\regs[30][0] ),
    .A1(\regs[31][0] ),
    .S(_02301_),
    .X(_03107_));
 sky130_fd_sc_hd__and2_1 _08700_ (.A(_02297_),
    .B(_03107_),
    .X(_03108_));
 sky130_fd_sc_hd__a211o_1 _08701_ (.A1(_02394_),
    .A2(_03106_),
    .B1(_03108_),
    .C1(_02538_),
    .X(_03109_));
 sky130_fd_sc_hd__or2b_1 _08702_ (.A(\regs[27][0] ),
    .B_N(_02333_),
    .X(_03110_));
 sky130_fd_sc_hd__o21a_1 _08703_ (.A1(_02333_),
    .A2(\regs[26][0] ),
    .B1(_02367_),
    .X(_03111_));
 sky130_fd_sc_hd__mux2_1 _08704_ (.A0(\regs[24][0] ),
    .A1(\regs[25][0] ),
    .S(_02458_),
    .X(_03112_));
 sky130_fd_sc_hd__a221o_1 _08705_ (.A1(_03110_),
    .A2(_03111_),
    .B1(_03112_),
    .B2(_02388_),
    .C1(_02293_),
    .X(_03113_));
 sky130_fd_sc_hd__a31o_1 _08706_ (.A1(_02290_),
    .A2(_03109_),
    .A3(_03113_),
    .B1(_02285_),
    .X(_03114_));
 sky130_fd_sc_hd__a21oi_1 _08707_ (.A1(_02365_),
    .A2(_03105_),
    .B1(_03114_),
    .Y(_03115_));
 sky130_fd_sc_hd__mux4_1 _08708_ (.A0(\regs[12][0] ),
    .A1(\regs[13][0] ),
    .A2(\regs[14][0] ),
    .A3(\regs[15][0] ),
    .S0(_02458_),
    .S1(_02297_),
    .X(_03116_));
 sky130_fd_sc_hd__or2_1 _08709_ (.A(_02330_),
    .B(_03116_),
    .X(_03117_));
 sky130_fd_sc_hd__mux4_1 _08710_ (.A0(\regs[8][0] ),
    .A1(\regs[9][0] ),
    .A2(\regs[10][0] ),
    .A3(\regs[11][0] ),
    .S0(_02354_),
    .S1(_02297_),
    .X(_03118_));
 sky130_fd_sc_hd__o21a_1 _08711_ (.A1(_02358_),
    .A2(_03118_),
    .B1(_02289_),
    .X(_03119_));
 sky130_fd_sc_hd__mux4_1 _08712_ (.A0(\regs[0][0] ),
    .A1(\regs[1][0] ),
    .A2(\regs[2][0] ),
    .A3(\regs[3][0] ),
    .S0(_02406_),
    .S1(_02297_),
    .X(_03120_));
 sky130_fd_sc_hd__mux4_1 _08713_ (.A0(\regs[4][0] ),
    .A1(\regs[5][0] ),
    .A2(\regs[6][0] ),
    .A3(\regs[7][0] ),
    .S0(_02406_),
    .S1(_02297_),
    .X(_03121_));
 sky130_fd_sc_hd__mux2_1 _08714_ (.A0(_03120_),
    .A1(_03121_),
    .S(_02358_),
    .X(_03122_));
 sky130_fd_sc_hd__a221o_1 _08715_ (.A1(_03117_),
    .A2(_03119_),
    .B1(_03122_),
    .B2(_02362_),
    .C1(_02433_),
    .X(_03123_));
 sky130_fd_sc_hd__or3b_2 _08716_ (.A(_02543_),
    .B(_03115_),
    .C_N(_03123_),
    .X(_03124_));
 sky130_fd_sc_hd__o21ai_1 _08717_ (.A1(_01776_),
    .A2(_00001_),
    .B1(_03124_),
    .Y(_01408_));
 sky130_fd_sc_hd__nor3b_4 _08718_ (.A(net1),
    .B(net34),
    .C_N(\core_state[3] ),
    .Y(_00000_));
 sky130_fd_sc_hd__inv_2 _08719_ (.A(\instret[50] ),
    .Y(_03125_));
 sky130_fd_sc_hd__inv_2 _08720_ (.A(\instret[49] ),
    .Y(_03126_));
 sky130_fd_sc_hd__inv_2 _08721_ (.A(\instret[48] ),
    .Y(_03127_));
 sky130_fd_sc_hd__and3_1 _08722_ (.A(\instret[2] ),
    .B(\instret[1] ),
    .C(\instret[0] ),
    .X(_03128_));
 sky130_fd_sc_hd__and2_1 _08723_ (.A(\instret[5] ),
    .B(\instret[4] ),
    .X(_03129_));
 sky130_fd_sc_hd__and4_1 _08724_ (.A(\instret[3] ),
    .B(_00000_),
    .C(_03128_),
    .D(_03129_),
    .X(_03130_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _08725_ (.A(_03130_),
    .X(_03131_));
 sky130_fd_sc_hd__and2_1 _08726_ (.A(\instret[7] ),
    .B(\instret[6] ),
    .X(_03132_));
 sky130_fd_sc_hd__and4_1 _08727_ (.A(\instret[9] ),
    .B(\instret[8] ),
    .C(_03131_),
    .D(_03132_),
    .X(_03133_));
 sky130_fd_sc_hd__and2_1 _08728_ (.A(\instret[13] ),
    .B(\instret[12] ),
    .X(_03134_));
 sky130_fd_sc_hd__and4_1 _08729_ (.A(\instret[11] ),
    .B(\instret[10] ),
    .C(_03133_),
    .D(_03134_),
    .X(_03135_));
 sky130_fd_sc_hd__and2_1 _08730_ (.A(\instret[15] ),
    .B(\instret[14] ),
    .X(_03136_));
 sky130_fd_sc_hd__and4_1 _08731_ (.A(\instret[17] ),
    .B(\instret[16] ),
    .C(_03135_),
    .D(_03136_),
    .X(_03137_));
 sky130_fd_sc_hd__and4_1 _08732_ (.A(\instret[20] ),
    .B(\instret[19] ),
    .C(\instret[18] ),
    .D(_03137_),
    .X(_03138_));
 sky130_fd_sc_hd__and4_1 _08733_ (.A(\instret[23] ),
    .B(\instret[22] ),
    .C(\instret[21] ),
    .D(_03138_),
    .X(_03139_));
 sky130_fd_sc_hd__and4_1 _08734_ (.A(\instret[26] ),
    .B(\instret[25] ),
    .C(\instret[24] ),
    .D(_03139_),
    .X(_03140_));
 sky130_fd_sc_hd__and4_1 _08735_ (.A(\instret[29] ),
    .B(\instret[28] ),
    .C(\instret[27] ),
    .D(_03140_),
    .X(_03141_));
 sky130_fd_sc_hd__and4_1 _08736_ (.A(\instret[32] ),
    .B(\instret[31] ),
    .C(\instret[30] ),
    .D(_03141_),
    .X(_03142_));
 sky130_fd_sc_hd__and4_2 _08737_ (.A(\instret[35] ),
    .B(\instret[34] ),
    .C(\instret[33] ),
    .D(_03142_),
    .X(_03143_));
 sky130_fd_sc_hd__and2_1 _08738_ (.A(\instret[37] ),
    .B(\instret[36] ),
    .X(_03144_));
 sky130_fd_sc_hd__and2_1 _08739_ (.A(\instret[39] ),
    .B(\instret[38] ),
    .X(_03145_));
 sky130_fd_sc_hd__and2_1 _08740_ (.A(\instret[41] ),
    .B(\instret[40] ),
    .X(_03146_));
 sky130_fd_sc_hd__and4_1 _08741_ (.A(_03143_),
    .B(_03144_),
    .C(_03145_),
    .D(_03146_),
    .X(_03147_));
 sky130_fd_sc_hd__buf_2 _08742_ (.A(_03147_),
    .X(_03148_));
 sky130_fd_sc_hd__and2_1 _08743_ (.A(\instret[43] ),
    .B(\instret[42] ),
    .X(_03149_));
 sky130_fd_sc_hd__and2_1 _08744_ (.A(\instret[45] ),
    .B(\instret[44] ),
    .X(_03150_));
 sky130_fd_sc_hd__and2_1 _08745_ (.A(\instret[47] ),
    .B(\instret[46] ),
    .X(_03151_));
 sky130_fd_sc_hd__nand4_4 _08746_ (.A(_03148_),
    .B(_03149_),
    .C(_03150_),
    .D(_03151_),
    .Y(_03152_));
 sky130_fd_sc_hd__nor4_2 _08747_ (.A(_03125_),
    .B(_03126_),
    .C(_03127_),
    .D(_03152_),
    .Y(_03153_));
 sky130_fd_sc_hd__and4_1 _08748_ (.A(\instret[53] ),
    .B(\instret[52] ),
    .C(\instret[51] ),
    .D(_03153_),
    .X(_03154_));
 sky130_fd_sc_hd__and4_1 _08749_ (.A(\instret[56] ),
    .B(\instret[55] ),
    .C(\instret[54] ),
    .D(_03154_),
    .X(_03155_));
 sky130_fd_sc_hd__and4_1 _08750_ (.A(\instret[59] ),
    .B(\instret[58] ),
    .C(\instret[57] ),
    .D(_03155_),
    .X(_03156_));
 sky130_fd_sc_hd__and4_1 _08751_ (.A(\instret[62] ),
    .B(\instret[61] ),
    .C(\instret[60] ),
    .D(_03156_),
    .X(_03157_));
 sky130_fd_sc_hd__xor2_1 _08752_ (.A(\instret[63] ),
    .B(_03157_),
    .X(_01407_));
 sky130_fd_sc_hd__and3_1 _08753_ (.A(\instret[61] ),
    .B(\instret[60] ),
    .C(_03156_),
    .X(_03158_));
 sky130_fd_sc_hd__xor2_1 _08754_ (.A(\instret[62] ),
    .B(_03158_),
    .X(_01406_));
 sky130_fd_sc_hd__a21oi_1 _08755_ (.A1(\instret[60] ),
    .A2(_03156_),
    .B1(\instret[61] ),
    .Y(_03159_));
 sky130_fd_sc_hd__nor2_1 _08756_ (.A(_03158_),
    .B(_03159_),
    .Y(_01405_));
 sky130_fd_sc_hd__xor2_1 _08757_ (.A(\instret[60] ),
    .B(_03156_),
    .X(_01404_));
 sky130_fd_sc_hd__a31o_1 _08758_ (.A1(\instret[58] ),
    .A2(\instret[57] ),
    .A3(_03155_),
    .B1(\instret[59] ),
    .X(_03160_));
 sky130_fd_sc_hd__and2b_1 _08759_ (.A_N(_03156_),
    .B(_03160_),
    .X(_03161_));
 sky130_fd_sc_hd__clkbuf_1 _08760_ (.A(_03161_),
    .X(_01403_));
 sky130_fd_sc_hd__nand2_1 _08761_ (.A(\instret[57] ),
    .B(_03155_),
    .Y(_03162_));
 sky130_fd_sc_hd__xnor2_1 _08762_ (.A(\instret[58] ),
    .B(_03162_),
    .Y(_01402_));
 sky130_fd_sc_hd__xor2_1 _08763_ (.A(\instret[57] ),
    .B(_03155_),
    .X(_01401_));
 sky130_fd_sc_hd__and3_1 _08764_ (.A(\instret[55] ),
    .B(\instret[54] ),
    .C(_03154_),
    .X(_03163_));
 sky130_fd_sc_hd__xor2_1 _08765_ (.A(\instret[56] ),
    .B(_03163_),
    .X(_01400_));
 sky130_fd_sc_hd__a21oi_1 _08766_ (.A1(\instret[54] ),
    .A2(_03154_),
    .B1(\instret[55] ),
    .Y(_03164_));
 sky130_fd_sc_hd__nor2_1 _08767_ (.A(_03163_),
    .B(_03164_),
    .Y(_01399_));
 sky130_fd_sc_hd__xor2_1 _08768_ (.A(\instret[54] ),
    .B(_03154_),
    .X(_01398_));
 sky130_fd_sc_hd__and3_1 _08769_ (.A(\instret[52] ),
    .B(\instret[51] ),
    .C(_03153_),
    .X(_03165_));
 sky130_fd_sc_hd__xor2_1 _08770_ (.A(\instret[53] ),
    .B(_03165_),
    .X(_01397_));
 sky130_fd_sc_hd__a21oi_1 _08771_ (.A1(\instret[51] ),
    .A2(_03153_),
    .B1(\instret[52] ),
    .Y(_03166_));
 sky130_fd_sc_hd__nor2_1 _08772_ (.A(_03165_),
    .B(_03166_),
    .Y(_01396_));
 sky130_fd_sc_hd__xor2_1 _08773_ (.A(\instret[51] ),
    .B(_03153_),
    .X(_01395_));
 sky130_fd_sc_hd__nor2_1 _08774_ (.A(_03127_),
    .B(_03152_),
    .Y(_03167_));
 sky130_fd_sc_hd__and2_1 _08775_ (.A(\instret[49] ),
    .B(_03167_),
    .X(_03168_));
 sky130_fd_sc_hd__nor2_1 _08776_ (.A(\instret[50] ),
    .B(_03168_),
    .Y(_03169_));
 sky130_fd_sc_hd__nor2_1 _08777_ (.A(_03153_),
    .B(_03169_),
    .Y(_01394_));
 sky130_fd_sc_hd__nor2_1 _08778_ (.A(\instret[49] ),
    .B(_03167_),
    .Y(_03170_));
 sky130_fd_sc_hd__nor2_1 _08779_ (.A(_03168_),
    .B(_03170_),
    .Y(_01393_));
 sky130_fd_sc_hd__xnor2_1 _08780_ (.A(\instret[48] ),
    .B(_03152_),
    .Y(_01392_));
 sky130_fd_sc_hd__and3_1 _08781_ (.A(_03148_),
    .B(_03149_),
    .C(_03150_),
    .X(_03171_));
 sky130_fd_sc_hd__and2_1 _08782_ (.A(\instret[46] ),
    .B(_03171_),
    .X(_03172_));
 sky130_fd_sc_hd__o21a_1 _08783_ (.A1(\instret[47] ),
    .A2(_03172_),
    .B1(_03152_),
    .X(_01391_));
 sky130_fd_sc_hd__nor2_1 _08784_ (.A(\instret[46] ),
    .B(_03171_),
    .Y(_03173_));
 sky130_fd_sc_hd__nor2_1 _08785_ (.A(_03172_),
    .B(_03173_),
    .Y(_01390_));
 sky130_fd_sc_hd__and2_1 _08786_ (.A(_03148_),
    .B(_03149_),
    .X(_03174_));
 sky130_fd_sc_hd__a21oi_1 _08787_ (.A1(\instret[44] ),
    .A2(_03174_),
    .B1(\instret[45] ),
    .Y(_03175_));
 sky130_fd_sc_hd__nor2_1 _08788_ (.A(_03171_),
    .B(_03175_),
    .Y(_01389_));
 sky130_fd_sc_hd__xor2_1 _08789_ (.A(\instret[44] ),
    .B(_03174_),
    .X(_01388_));
 sky130_fd_sc_hd__a21oi_1 _08790_ (.A1(\instret[42] ),
    .A2(_03148_),
    .B1(\instret[43] ),
    .Y(_03176_));
 sky130_fd_sc_hd__nor2_1 _08791_ (.A(_03174_),
    .B(_03176_),
    .Y(_01387_));
 sky130_fd_sc_hd__xor2_1 _08792_ (.A(\instret[42] ),
    .B(_03148_),
    .X(_01386_));
 sky130_fd_sc_hd__and3_1 _08793_ (.A(_03143_),
    .B(_03144_),
    .C(_03145_),
    .X(_03177_));
 sky130_fd_sc_hd__and2_1 _08794_ (.A(\instret[40] ),
    .B(_03177_),
    .X(_03178_));
 sky130_fd_sc_hd__o21ba_1 _08795_ (.A1(\instret[41] ),
    .A2(_03178_),
    .B1_N(_03148_),
    .X(_01385_));
 sky130_fd_sc_hd__nor2_1 _08796_ (.A(\instret[40] ),
    .B(_03177_),
    .Y(_03179_));
 sky130_fd_sc_hd__nor2_1 _08797_ (.A(_03178_),
    .B(_03179_),
    .Y(_01384_));
 sky130_fd_sc_hd__and3_1 _08798_ (.A(\instret[38] ),
    .B(_03143_),
    .C(_03144_),
    .X(_03180_));
 sky130_fd_sc_hd__o21ba_1 _08799_ (.A1(\instret[39] ),
    .A2(_03180_),
    .B1_N(_03177_),
    .X(_01383_));
 sky130_fd_sc_hd__and2_1 _08800_ (.A(_03143_),
    .B(_03144_),
    .X(_03181_));
 sky130_fd_sc_hd__nor2_1 _08801_ (.A(\instret[38] ),
    .B(_03181_),
    .Y(_03182_));
 sky130_fd_sc_hd__nor2_1 _08802_ (.A(_03180_),
    .B(_03182_),
    .Y(_01382_));
 sky130_fd_sc_hd__a21oi_1 _08803_ (.A1(\instret[36] ),
    .A2(_03143_),
    .B1(\instret[37] ),
    .Y(_03183_));
 sky130_fd_sc_hd__nor2_1 _08804_ (.A(_03181_),
    .B(_03183_),
    .Y(_01381_));
 sky130_fd_sc_hd__xor2_1 _08805_ (.A(\instret[36] ),
    .B(_03143_),
    .X(_01380_));
 sky130_fd_sc_hd__a31o_1 _08806_ (.A1(\instret[34] ),
    .A2(\instret[33] ),
    .A3(_03142_),
    .B1(\instret[35] ),
    .X(_03184_));
 sky130_fd_sc_hd__and2b_1 _08807_ (.A_N(_03143_),
    .B(_03184_),
    .X(_03185_));
 sky130_fd_sc_hd__clkbuf_1 _08808_ (.A(_03185_),
    .X(_01379_));
 sky130_fd_sc_hd__nand2_1 _08809_ (.A(\instret[33] ),
    .B(_03142_),
    .Y(_03186_));
 sky130_fd_sc_hd__xnor2_1 _08810_ (.A(\instret[34] ),
    .B(_03186_),
    .Y(_01378_));
 sky130_fd_sc_hd__or2_1 _08811_ (.A(\instret[33] ),
    .B(_03142_),
    .X(_03187_));
 sky130_fd_sc_hd__and2_1 _08812_ (.A(_03186_),
    .B(_03187_),
    .X(_03188_));
 sky130_fd_sc_hd__clkbuf_1 _08813_ (.A(_03188_),
    .X(_01377_));
 sky130_fd_sc_hd__a31o_1 _08814_ (.A1(\instret[31] ),
    .A2(\instret[30] ),
    .A3(_03141_),
    .B1(\instret[32] ),
    .X(_03189_));
 sky130_fd_sc_hd__and2b_1 _08815_ (.A_N(_03142_),
    .B(_03189_),
    .X(_03190_));
 sky130_fd_sc_hd__clkbuf_1 _08816_ (.A(_03190_),
    .X(_01376_));
 sky130_fd_sc_hd__nand2_1 _08817_ (.A(\instret[30] ),
    .B(_03141_),
    .Y(_03191_));
 sky130_fd_sc_hd__xnor2_1 _08818_ (.A(\instret[31] ),
    .B(_03191_),
    .Y(_01375_));
 sky130_fd_sc_hd__or2_1 _08819_ (.A(\instret[30] ),
    .B(_03141_),
    .X(_03192_));
 sky130_fd_sc_hd__and2_1 _08820_ (.A(_03191_),
    .B(_03192_),
    .X(_03193_));
 sky130_fd_sc_hd__clkbuf_1 _08821_ (.A(_03193_),
    .X(_01374_));
 sky130_fd_sc_hd__a31o_1 _08822_ (.A1(\instret[28] ),
    .A2(\instret[27] ),
    .A3(_03140_),
    .B1(\instret[29] ),
    .X(_03194_));
 sky130_fd_sc_hd__and2b_1 _08823_ (.A_N(_03141_),
    .B(_03194_),
    .X(_03195_));
 sky130_fd_sc_hd__clkbuf_1 _08824_ (.A(_03195_),
    .X(_01373_));
 sky130_fd_sc_hd__nand2_1 _08825_ (.A(\instret[27] ),
    .B(_03140_),
    .Y(_03196_));
 sky130_fd_sc_hd__xnor2_1 _08826_ (.A(\instret[28] ),
    .B(_03196_),
    .Y(_01372_));
 sky130_fd_sc_hd__or2_1 _08827_ (.A(\instret[27] ),
    .B(_03140_),
    .X(_03197_));
 sky130_fd_sc_hd__and2_1 _08828_ (.A(_03196_),
    .B(_03197_),
    .X(_03198_));
 sky130_fd_sc_hd__clkbuf_1 _08829_ (.A(_03198_),
    .X(_01371_));
 sky130_fd_sc_hd__a31o_1 _08830_ (.A1(\instret[25] ),
    .A2(\instret[24] ),
    .A3(_03139_),
    .B1(\instret[26] ),
    .X(_03199_));
 sky130_fd_sc_hd__and2b_1 _08831_ (.A_N(_03140_),
    .B(_03199_),
    .X(_03200_));
 sky130_fd_sc_hd__clkbuf_1 _08832_ (.A(_03200_),
    .X(_01370_));
 sky130_fd_sc_hd__and2_1 _08833_ (.A(\instret[24] ),
    .B(_03139_),
    .X(_03201_));
 sky130_fd_sc_hd__xor2_1 _08834_ (.A(\instret[25] ),
    .B(_03201_),
    .X(_01369_));
 sky130_fd_sc_hd__nor2_1 _08835_ (.A(\instret[24] ),
    .B(_03139_),
    .Y(_03202_));
 sky130_fd_sc_hd__nor2_1 _08836_ (.A(_03201_),
    .B(_03202_),
    .Y(_01368_));
 sky130_fd_sc_hd__and3_1 _08837_ (.A(\instret[22] ),
    .B(\instret[21] ),
    .C(_03138_),
    .X(_03203_));
 sky130_fd_sc_hd__nor2_1 _08838_ (.A(\instret[23] ),
    .B(_03203_),
    .Y(_03204_));
 sky130_fd_sc_hd__nor2_1 _08839_ (.A(_03139_),
    .B(_03204_),
    .Y(_01367_));
 sky130_fd_sc_hd__a21oi_1 _08840_ (.A1(\instret[21] ),
    .A2(_03138_),
    .B1(\instret[22] ),
    .Y(_03205_));
 sky130_fd_sc_hd__nor2_1 _08841_ (.A(_03203_),
    .B(_03205_),
    .Y(_01366_));
 sky130_fd_sc_hd__xor2_1 _08842_ (.A(\instret[21] ),
    .B(_03138_),
    .X(_01365_));
 sky130_fd_sc_hd__a31o_1 _08843_ (.A1(\instret[19] ),
    .A2(\instret[18] ),
    .A3(_03137_),
    .B1(\instret[20] ),
    .X(_03206_));
 sky130_fd_sc_hd__and2b_1 _08844_ (.A_N(_03138_),
    .B(_03206_),
    .X(_03207_));
 sky130_fd_sc_hd__clkbuf_1 _08845_ (.A(_03207_),
    .X(_01364_));
 sky130_fd_sc_hd__nand2_1 _08846_ (.A(\instret[18] ),
    .B(_03137_),
    .Y(_03208_));
 sky130_fd_sc_hd__xnor2_1 _08847_ (.A(\instret[19] ),
    .B(_03208_),
    .Y(_01363_));
 sky130_fd_sc_hd__or2_1 _08848_ (.A(\instret[18] ),
    .B(_03137_),
    .X(_03209_));
 sky130_fd_sc_hd__and2_1 _08849_ (.A(_03208_),
    .B(_03209_),
    .X(_03210_));
 sky130_fd_sc_hd__clkbuf_1 _08850_ (.A(_03210_),
    .X(_01362_));
 sky130_fd_sc_hd__a31o_1 _08851_ (.A1(\instret[16] ),
    .A2(_03135_),
    .A3(_03136_),
    .B1(\instret[17] ),
    .X(_03211_));
 sky130_fd_sc_hd__and2b_1 _08852_ (.A_N(_03137_),
    .B(_03211_),
    .X(_03212_));
 sky130_fd_sc_hd__clkbuf_1 _08853_ (.A(_03212_),
    .X(_01361_));
 sky130_fd_sc_hd__nand2_1 _08854_ (.A(_03135_),
    .B(_03136_),
    .Y(_03213_));
 sky130_fd_sc_hd__xnor2_1 _08855_ (.A(\instret[16] ),
    .B(_03213_),
    .Y(_01360_));
 sky130_fd_sc_hd__a21o_1 _08856_ (.A1(\instret[14] ),
    .A2(_03135_),
    .B1(\instret[15] ),
    .X(_03214_));
 sky130_fd_sc_hd__and2_1 _08857_ (.A(_03213_),
    .B(_03214_),
    .X(_03215_));
 sky130_fd_sc_hd__clkbuf_1 _08858_ (.A(_03215_),
    .X(_01359_));
 sky130_fd_sc_hd__xor2_1 _08859_ (.A(\instret[14] ),
    .B(_03135_),
    .X(_01358_));
 sky130_fd_sc_hd__and3_1 _08860_ (.A(\instret[11] ),
    .B(\instret[10] ),
    .C(_03133_),
    .X(_03216_));
 sky130_fd_sc_hd__and2_1 _08861_ (.A(\instret[12] ),
    .B(_03216_),
    .X(_03217_));
 sky130_fd_sc_hd__o21ba_1 _08862_ (.A1(\instret[13] ),
    .A2(_03217_),
    .B1_N(_03135_),
    .X(_01357_));
 sky130_fd_sc_hd__nor2_1 _08863_ (.A(\instret[12] ),
    .B(_03216_),
    .Y(_03218_));
 sky130_fd_sc_hd__nor2_1 _08864_ (.A(_03217_),
    .B(_03218_),
    .Y(_01356_));
 sky130_fd_sc_hd__a21oi_1 _08865_ (.A1(\instret[10] ),
    .A2(_03133_),
    .B1(\instret[11] ),
    .Y(_03219_));
 sky130_fd_sc_hd__nor2_1 _08866_ (.A(_03216_),
    .B(_03219_),
    .Y(_01355_));
 sky130_fd_sc_hd__xor2_1 _08867_ (.A(\instret[10] ),
    .B(_03133_),
    .X(_01354_));
 sky130_fd_sc_hd__a31o_1 _08868_ (.A1(\instret[8] ),
    .A2(_03131_),
    .A3(_03132_),
    .B1(\instret[9] ),
    .X(_03220_));
 sky130_fd_sc_hd__and2b_1 _08869_ (.A_N(_03133_),
    .B(_03220_),
    .X(_03221_));
 sky130_fd_sc_hd__clkbuf_1 _08870_ (.A(_03221_),
    .X(_01353_));
 sky130_fd_sc_hd__and2_1 _08871_ (.A(_03131_),
    .B(_03132_),
    .X(_03222_));
 sky130_fd_sc_hd__xor2_1 _08872_ (.A(\instret[8] ),
    .B(_03222_),
    .X(_01352_));
 sky130_fd_sc_hd__a21oi_1 _08873_ (.A1(\instret[6] ),
    .A2(_03131_),
    .B1(\instret[7] ),
    .Y(_03223_));
 sky130_fd_sc_hd__nor2_1 _08874_ (.A(_03222_),
    .B(_03223_),
    .Y(_01351_));
 sky130_fd_sc_hd__xor2_1 _08875_ (.A(\instret[6] ),
    .B(_03131_),
    .X(_01350_));
 sky130_fd_sc_hd__and3_1 _08876_ (.A(\instret[3] ),
    .B(_00000_),
    .C(_03128_),
    .X(_03224_));
 sky130_fd_sc_hd__and2_1 _08877_ (.A(\instret[4] ),
    .B(_03224_),
    .X(_03225_));
 sky130_fd_sc_hd__o21ba_1 _08878_ (.A1(\instret[5] ),
    .A2(_03225_),
    .B1_N(_03131_),
    .X(_01349_));
 sky130_fd_sc_hd__nor2_1 _08879_ (.A(\instret[4] ),
    .B(_03224_),
    .Y(_03226_));
 sky130_fd_sc_hd__nor2_1 _08880_ (.A(_03225_),
    .B(_03226_),
    .Y(_01348_));
 sky130_fd_sc_hd__a21oi_1 _08881_ (.A1(_00000_),
    .A2(_03128_),
    .B1(\instret[3] ),
    .Y(_03227_));
 sky130_fd_sc_hd__nor2_1 _08882_ (.A(_03224_),
    .B(_03227_),
    .Y(_01347_));
 sky130_fd_sc_hd__and3_1 _08883_ (.A(\instret[1] ),
    .B(\instret[0] ),
    .C(_00000_),
    .X(_03228_));
 sky130_fd_sc_hd__o2bb2a_1 _08884_ (.A1_N(_00000_),
    .A2_N(_03128_),
    .B1(_03228_),
    .B2(\instret[2] ),
    .X(_01346_));
 sky130_fd_sc_hd__a21oi_1 _08885_ (.A1(\instret[0] ),
    .A2(_00000_),
    .B1(\instret[1] ),
    .Y(_03229_));
 sky130_fd_sc_hd__nor2_1 _08886_ (.A(_03228_),
    .B(_03229_),
    .Y(_01345_));
 sky130_fd_sc_hd__nand2_1 _08887_ (.A(\instret[0] ),
    .B(_00000_),
    .Y(_03230_));
 sky130_fd_sc_hd__or2_1 _08888_ (.A(\instret[0] ),
    .B(_00000_),
    .X(_03231_));
 sky130_fd_sc_hd__and2_1 _08889_ (.A(_03230_),
    .B(_03231_),
    .X(_03232_));
 sky130_fd_sc_hd__clkbuf_1 _08890_ (.A(_03232_),
    .X(_01344_));
 sky130_fd_sc_hd__buf_6 _08891_ (.A(net18),
    .X(_03233_));
 sky130_fd_sc_hd__inv_2 _08892_ (.A(net16),
    .Y(_03234_));
 sky130_fd_sc_hd__buf_6 _08893_ (.A(_03234_),
    .X(_03235_));
 sky130_fd_sc_hd__buf_8 _08894_ (.A(_03235_),
    .X(_03236_));
 sky130_fd_sc_hd__buf_8 _08895_ (.A(net14),
    .X(_03237_));
 sky130_fd_sc_hd__buf_8 _08896_ (.A(_03237_),
    .X(_03238_));
 sky130_fd_sc_hd__buf_8 _08897_ (.A(net15),
    .X(_03239_));
 sky130_fd_sc_hd__buf_6 _08898_ (.A(_03239_),
    .X(_03240_));
 sky130_fd_sc_hd__mux4_1 _08899_ (.A0(\regs[12][31] ),
    .A1(\regs[13][31] ),
    .A2(\regs[14][31] ),
    .A3(\regs[15][31] ),
    .S0(_03238_),
    .S1(_03240_),
    .X(_03241_));
 sky130_fd_sc_hd__or2_1 _08900_ (.A(_03236_),
    .B(_03241_),
    .X(_03242_));
 sky130_fd_sc_hd__buf_6 _08901_ (.A(net16),
    .X(_03243_));
 sky130_fd_sc_hd__clkbuf_8 _08902_ (.A(_03243_),
    .X(_03244_));
 sky130_fd_sc_hd__buf_6 _08903_ (.A(net15),
    .X(_03245_));
 sky130_fd_sc_hd__buf_6 _08904_ (.A(_03245_),
    .X(_03246_));
 sky130_fd_sc_hd__mux4_1 _08905_ (.A0(\regs[8][31] ),
    .A1(\regs[9][31] ),
    .A2(\regs[10][31] ),
    .A3(\regs[11][31] ),
    .S0(_03238_),
    .S1(_03246_),
    .X(_03247_));
 sky130_fd_sc_hd__o21a_1 _08906_ (.A1(_03244_),
    .A2(_03247_),
    .B1(_02267_),
    .X(_03248_));
 sky130_fd_sc_hd__buf_8 _08907_ (.A(_03237_),
    .X(_03249_));
 sky130_fd_sc_hd__buf_6 _08908_ (.A(net15),
    .X(_03250_));
 sky130_fd_sc_hd__buf_8 _08909_ (.A(_03250_),
    .X(_03251_));
 sky130_fd_sc_hd__mux4_1 _08910_ (.A0(\regs[0][31] ),
    .A1(\regs[1][31] ),
    .A2(\regs[2][31] ),
    .A3(\regs[3][31] ),
    .S0(_03249_),
    .S1(_03251_),
    .X(_03252_));
 sky130_fd_sc_hd__mux4_1 _08911_ (.A0(\regs[4][31] ),
    .A1(\regs[5][31] ),
    .A2(\regs[6][31] ),
    .A3(\regs[7][31] ),
    .S0(_03249_),
    .S1(_03251_),
    .X(_03253_));
 sky130_fd_sc_hd__buf_6 _08912_ (.A(net16),
    .X(_03254_));
 sky130_fd_sc_hd__buf_6 _08913_ (.A(_03254_),
    .X(_03255_));
 sky130_fd_sc_hd__mux2_1 _08914_ (.A0(_03252_),
    .A1(_03253_),
    .S(_03255_),
    .X(_03256_));
 sky130_fd_sc_hd__inv_2 _08915_ (.A(net17),
    .Y(_03257_));
 sky130_fd_sc_hd__buf_6 _08916_ (.A(_03257_),
    .X(_03258_));
 sky130_fd_sc_hd__buf_6 _08917_ (.A(_03258_),
    .X(_03259_));
 sky130_fd_sc_hd__a22o_1 _08918_ (.A1(_03242_),
    .A2(_03248_),
    .B1(_03256_),
    .B2(_03259_),
    .X(_03260_));
 sky130_fd_sc_hd__buf_8 _08919_ (.A(_02281_),
    .X(_03261_));
 sky130_fd_sc_hd__buf_8 _08920_ (.A(_02276_),
    .X(_03262_));
 sky130_fd_sc_hd__mux4_1 _08921_ (.A0(\regs[16][31] ),
    .A1(\regs[17][31] ),
    .A2(\regs[18][31] ),
    .A3(\regs[19][31] ),
    .S0(_03261_),
    .S1(_03262_),
    .X(_03263_));
 sky130_fd_sc_hd__mux4_1 _08922_ (.A0(\regs[20][31] ),
    .A1(\regs[21][31] ),
    .A2(\regs[22][31] ),
    .A3(\regs[23][31] ),
    .S0(_02282_),
    .S1(_03262_),
    .X(_03264_));
 sky130_fd_sc_hd__mux2_1 _08923_ (.A0(_03263_),
    .A1(_03264_),
    .S(_02272_),
    .X(_03265_));
 sky130_fd_sc_hd__clkbuf_8 _08924_ (.A(net17),
    .X(_03266_));
 sky130_fd_sc_hd__buf_6 _08925_ (.A(_03266_),
    .X(_03267_));
 sky130_fd_sc_hd__clkbuf_16 _08926_ (.A(_02276_),
    .X(_03268_));
 sky130_fd_sc_hd__buf_6 _08927_ (.A(net14),
    .X(_03269_));
 sky130_fd_sc_hd__buf_6 _08928_ (.A(_03269_),
    .X(_03270_));
 sky130_fd_sc_hd__mux2_1 _08929_ (.A0(\regs[30][31] ),
    .A1(\regs[31][31] ),
    .S(_03270_),
    .X(_03271_));
 sky130_fd_sc_hd__inv_4 _08930_ (.A(net15),
    .Y(_03272_));
 sky130_fd_sc_hd__mux2_1 _08931_ (.A0(\regs[28][31] ),
    .A1(\regs[29][31] ),
    .S(_03269_),
    .X(_03273_));
 sky130_fd_sc_hd__clkbuf_8 _08932_ (.A(_03234_),
    .X(_03274_));
 sky130_fd_sc_hd__a21o_1 _08933_ (.A1(_03272_),
    .A2(_03273_),
    .B1(_03274_),
    .X(_03275_));
 sky130_fd_sc_hd__a21o_1 _08934_ (.A1(_03268_),
    .A2(_03271_),
    .B1(_03275_),
    .X(_03276_));
 sky130_fd_sc_hd__clkbuf_8 _08935_ (.A(_03237_),
    .X(_03277_));
 sky130_fd_sc_hd__or2b_1 _08936_ (.A(\regs[27][31] ),
    .B_N(_03277_),
    .X(_03278_));
 sky130_fd_sc_hd__o21a_1 _08937_ (.A1(_03277_),
    .A2(\regs[26][31] ),
    .B1(_02276_),
    .X(_03279_));
 sky130_fd_sc_hd__clkbuf_8 _08938_ (.A(_02280_),
    .X(_03280_));
 sky130_fd_sc_hd__mux2_1 _08939_ (.A0(\regs[24][31] ),
    .A1(\regs[25][31] ),
    .S(_03280_),
    .X(_03281_));
 sky130_fd_sc_hd__buf_4 _08940_ (.A(_03272_),
    .X(_03282_));
 sky130_fd_sc_hd__a221o_1 _08941_ (.A1(_03278_),
    .A2(_03279_),
    .B1(_03281_),
    .B2(_03282_),
    .C1(_03243_),
    .X(_03283_));
 sky130_fd_sc_hd__a31o_1 _08942_ (.A1(_03267_),
    .A2(_03276_),
    .A3(_03283_),
    .B1(_02263_),
    .X(_03284_));
 sky130_fd_sc_hd__a21o_1 _08943_ (.A1(_03259_),
    .A2(_03265_),
    .B1(_03284_),
    .X(_03285_));
 sky130_fd_sc_hd__o211a_1 _08944_ (.A1(_03233_),
    .A2(_03260_),
    .B1(_03285_),
    .C1(_02254_),
    .X(_03286_));
 sky130_fd_sc_hd__a21o_1 _08945_ (.A1(\rs2_content[31] ),
    .A2(_02543_),
    .B1(_03286_),
    .X(_01343_));
 sky130_fd_sc_hd__buf_6 _08946_ (.A(_03234_),
    .X(_03287_));
 sky130_fd_sc_hd__buf_6 _08947_ (.A(_03287_),
    .X(_03288_));
 sky130_fd_sc_hd__buf_6 _08948_ (.A(_03269_),
    .X(_03289_));
 sky130_fd_sc_hd__buf_6 _08949_ (.A(_03289_),
    .X(_03290_));
 sky130_fd_sc_hd__buf_8 _08950_ (.A(_03251_),
    .X(_03291_));
 sky130_fd_sc_hd__mux4_1 _08951_ (.A0(\regs[12][30] ),
    .A1(\regs[13][30] ),
    .A2(\regs[14][30] ),
    .A3(\regs[15][30] ),
    .S0(_03290_),
    .S1(_03291_),
    .X(_03292_));
 sky130_fd_sc_hd__or2_1 _08952_ (.A(_03288_),
    .B(_03292_),
    .X(_03293_));
 sky130_fd_sc_hd__clkbuf_16 _08953_ (.A(_03249_),
    .X(_03294_));
 sky130_fd_sc_hd__buf_8 _08954_ (.A(_03240_),
    .X(_03295_));
 sky130_fd_sc_hd__mux4_1 _08955_ (.A0(\regs[8][30] ),
    .A1(\regs[9][30] ),
    .A2(\regs[10][30] ),
    .A3(\regs[11][30] ),
    .S0(_03294_),
    .S1(_03295_),
    .X(_03296_));
 sky130_fd_sc_hd__buf_6 _08956_ (.A(_03266_),
    .X(_03297_));
 sky130_fd_sc_hd__o21a_1 _08957_ (.A1(_02273_),
    .A2(_03296_),
    .B1(_03297_),
    .X(_03298_));
 sky130_fd_sc_hd__buf_12 _08958_ (.A(_02280_),
    .X(_03299_));
 sky130_fd_sc_hd__clkbuf_16 _08959_ (.A(_03299_),
    .X(_03300_));
 sky130_fd_sc_hd__buf_8 _08960_ (.A(_03251_),
    .X(_03301_));
 sky130_fd_sc_hd__mux4_1 _08961_ (.A0(\regs[0][30] ),
    .A1(\regs[1][30] ),
    .A2(\regs[2][30] ),
    .A3(\regs[3][30] ),
    .S0(_03300_),
    .S1(_03301_),
    .X(_03302_));
 sky130_fd_sc_hd__clkbuf_16 _08962_ (.A(_03299_),
    .X(_03303_));
 sky130_fd_sc_hd__buf_6 _08963_ (.A(_03250_),
    .X(_03304_));
 sky130_fd_sc_hd__buf_8 _08964_ (.A(_03304_),
    .X(_03305_));
 sky130_fd_sc_hd__mux4_1 _08965_ (.A0(\regs[4][30] ),
    .A1(\regs[5][30] ),
    .A2(\regs[6][30] ),
    .A3(\regs[7][30] ),
    .S0(_03303_),
    .S1(_03305_),
    .X(_03306_));
 sky130_fd_sc_hd__buf_8 _08966_ (.A(_03243_),
    .X(_03307_));
 sky130_fd_sc_hd__mux2_1 _08967_ (.A0(_03302_),
    .A1(_03306_),
    .S(_03307_),
    .X(_03308_));
 sky130_fd_sc_hd__buf_6 _08968_ (.A(_03258_),
    .X(_03309_));
 sky130_fd_sc_hd__buf_6 _08969_ (.A(_03309_),
    .X(_03310_));
 sky130_fd_sc_hd__a22o_1 _08970_ (.A1(_03293_),
    .A2(_03298_),
    .B1(_03308_),
    .B2(_03310_),
    .X(_03311_));
 sky130_fd_sc_hd__clkbuf_8 _08971_ (.A(_03259_),
    .X(_03312_));
 sky130_fd_sc_hd__buf_6 _08972_ (.A(_03262_),
    .X(_03313_));
 sky130_fd_sc_hd__mux4_1 _08973_ (.A0(\regs[16][30] ),
    .A1(\regs[17][30] ),
    .A2(\regs[18][30] ),
    .A3(\regs[19][30] ),
    .S0(_02283_),
    .S1(_03313_),
    .X(_03314_));
 sky130_fd_sc_hd__mux4_1 _08974_ (.A0(\regs[20][30] ),
    .A1(\regs[21][30] ),
    .A2(\regs[22][30] ),
    .A3(\regs[23][30] ),
    .S0(_02283_),
    .S1(_03313_),
    .X(_03315_));
 sky130_fd_sc_hd__buf_6 _08975_ (.A(_02272_),
    .X(_03316_));
 sky130_fd_sc_hd__mux2_1 _08976_ (.A0(_03314_),
    .A1(_03315_),
    .S(_03316_),
    .X(_03317_));
 sky130_fd_sc_hd__buf_8 _08977_ (.A(_03299_),
    .X(_03318_));
 sky130_fd_sc_hd__mux2_1 _08978_ (.A0(\regs[30][30] ),
    .A1(\regs[31][30] ),
    .S(_03318_),
    .X(_03319_));
 sky130_fd_sc_hd__clkbuf_8 _08979_ (.A(_03272_),
    .X(_03320_));
 sky130_fd_sc_hd__mux2_1 _08980_ (.A0(\regs[28][30] ),
    .A1(\regs[29][30] ),
    .S(_03289_),
    .X(_03321_));
 sky130_fd_sc_hd__a21o_1 _08981_ (.A1(_03320_),
    .A2(_03321_),
    .B1(_03287_),
    .X(_03322_));
 sky130_fd_sc_hd__a21o_1 _08982_ (.A1(_02278_),
    .A2(_03319_),
    .B1(_03322_),
    .X(_03323_));
 sky130_fd_sc_hd__clkbuf_4 _08983_ (.A(_03277_),
    .X(_03324_));
 sky130_fd_sc_hd__or2b_1 _08984_ (.A(\regs[27][30] ),
    .B_N(_03324_),
    .X(_03325_));
 sky130_fd_sc_hd__o21a_1 _08985_ (.A1(_03290_),
    .A2(\regs[26][30] ),
    .B1(_02277_),
    .X(_03326_));
 sky130_fd_sc_hd__buf_6 _08986_ (.A(_03280_),
    .X(_03327_));
 sky130_fd_sc_hd__mux2_1 _08987_ (.A0(\regs[24][30] ),
    .A1(\regs[25][30] ),
    .S(_03327_),
    .X(_03328_));
 sky130_fd_sc_hd__buf_4 _08988_ (.A(_03282_),
    .X(_03329_));
 sky130_fd_sc_hd__a221o_1 _08989_ (.A1(_03325_),
    .A2(_03326_),
    .B1(_03328_),
    .B2(_03329_),
    .C1(_03244_),
    .X(_03330_));
 sky130_fd_sc_hd__nand2_4 _08990_ (.A(_03233_),
    .B(_02252_),
    .Y(_03331_));
 sky130_fd_sc_hd__a31o_1 _08991_ (.A1(_02268_),
    .A2(_03323_),
    .A3(_03330_),
    .B1(_03331_),
    .X(_03332_));
 sky130_fd_sc_hd__a21o_1 _08992_ (.A1(_03312_),
    .A2(_03317_),
    .B1(_03332_),
    .X(_03333_));
 sky130_fd_sc_hd__o221a_1 _08993_ (.A1(\rs2_content[30] ),
    .A2(_02754_),
    .B1(_02266_),
    .B2(_03311_),
    .C1(_03333_),
    .X(_01342_));
 sky130_fd_sc_hd__buf_6 _08994_ (.A(_03309_),
    .X(_03334_));
 sky130_fd_sc_hd__buf_8 _08995_ (.A(_03299_),
    .X(_03335_));
 sky130_fd_sc_hd__buf_6 _08996_ (.A(_03304_),
    .X(_03336_));
 sky130_fd_sc_hd__mux4_1 _08997_ (.A0(\regs[16][29] ),
    .A1(\regs[17][29] ),
    .A2(\regs[18][29] ),
    .A3(\regs[19][29] ),
    .S0(_03335_),
    .S1(_03336_),
    .X(_03337_));
 sky130_fd_sc_hd__mux4_1 _08998_ (.A0(\regs[20][29] ),
    .A1(\regs[21][29] ),
    .A2(\regs[22][29] ),
    .A3(\regs[23][29] ),
    .S0(_03335_),
    .S1(_03336_),
    .X(_03338_));
 sky130_fd_sc_hd__clkbuf_16 _08999_ (.A(_03243_),
    .X(_03339_));
 sky130_fd_sc_hd__mux2_1 _09000_ (.A0(_03337_),
    .A1(_03338_),
    .S(_03339_),
    .X(_03340_));
 sky130_fd_sc_hd__buf_6 _09001_ (.A(_03304_),
    .X(_03341_));
 sky130_fd_sc_hd__buf_6 _09002_ (.A(_02280_),
    .X(_03342_));
 sky130_fd_sc_hd__buf_4 _09003_ (.A(_03342_),
    .X(_03343_));
 sky130_fd_sc_hd__mux2_1 _09004_ (.A0(\regs[30][29] ),
    .A1(\regs[31][29] ),
    .S(_03343_),
    .X(_03344_));
 sky130_fd_sc_hd__and2_1 _09005_ (.A(_03341_),
    .B(_03344_),
    .X(_03345_));
 sky130_fd_sc_hd__buf_4 _09006_ (.A(_03342_),
    .X(_03346_));
 sky130_fd_sc_hd__mux2_1 _09007_ (.A0(\regs[28][29] ),
    .A1(\regs[29][29] ),
    .S(_03346_),
    .X(_03347_));
 sky130_fd_sc_hd__a21o_1 _09008_ (.A1(_03329_),
    .A2(_03347_),
    .B1(_03236_),
    .X(_03348_));
 sky130_fd_sc_hd__buf_6 _09009_ (.A(_02280_),
    .X(_03349_));
 sky130_fd_sc_hd__buf_4 _09010_ (.A(_03349_),
    .X(_03350_));
 sky130_fd_sc_hd__or2b_1 _09011_ (.A(\regs[27][29] ),
    .B_N(_03350_),
    .X(_03351_));
 sky130_fd_sc_hd__buf_6 _09012_ (.A(_03245_),
    .X(_03352_));
 sky130_fd_sc_hd__o21a_1 _09013_ (.A1(_03350_),
    .A2(\regs[26][29] ),
    .B1(_03352_),
    .X(_03353_));
 sky130_fd_sc_hd__mux2_1 _09014_ (.A0(\regs[24][29] ),
    .A1(\regs[25][29] ),
    .S(_03343_),
    .X(_03354_));
 sky130_fd_sc_hd__buf_4 _09015_ (.A(_03272_),
    .X(_03355_));
 sky130_fd_sc_hd__buf_4 _09016_ (.A(_03355_),
    .X(_03356_));
 sky130_fd_sc_hd__buf_6 _09017_ (.A(_02271_),
    .X(_03357_));
 sky130_fd_sc_hd__a221o_1 _09018_ (.A1(_03351_),
    .A2(_03353_),
    .B1(_03354_),
    .B2(_03356_),
    .C1(_03357_),
    .X(_03358_));
 sky130_fd_sc_hd__buf_6 _09019_ (.A(_02267_),
    .X(_03359_));
 sky130_fd_sc_hd__o211a_1 _09020_ (.A1(_03345_),
    .A2(_03348_),
    .B1(_03358_),
    .C1(_03359_),
    .X(_03360_));
 sky130_fd_sc_hd__a211o_1 _09021_ (.A1(_03334_),
    .A2(_03340_),
    .B1(_03360_),
    .C1(_02264_),
    .X(_03361_));
 sky130_fd_sc_hd__clkbuf_8 _09022_ (.A(_03287_),
    .X(_03362_));
 sky130_fd_sc_hd__buf_12 _09023_ (.A(_03299_),
    .X(_03363_));
 sky130_fd_sc_hd__mux4_1 _09024_ (.A0(\regs[12][29] ),
    .A1(\regs[13][29] ),
    .A2(\regs[14][29] ),
    .A3(\regs[15][29] ),
    .S0(_03363_),
    .S1(_03268_),
    .X(_03364_));
 sky130_fd_sc_hd__or2_1 _09025_ (.A(_03362_),
    .B(_03364_),
    .X(_03365_));
 sky130_fd_sc_hd__buf_6 _09026_ (.A(_03255_),
    .X(_03366_));
 sky130_fd_sc_hd__mux4_1 _09027_ (.A0(\regs[8][29] ),
    .A1(\regs[9][29] ),
    .A2(\regs[10][29] ),
    .A3(\regs[11][29] ),
    .S0(_03300_),
    .S1(_03301_),
    .X(_03367_));
 sky130_fd_sc_hd__clkbuf_8 _09028_ (.A(_03266_),
    .X(_03368_));
 sky130_fd_sc_hd__o21a_1 _09029_ (.A1(_03366_),
    .A2(_03367_),
    .B1(_03368_),
    .X(_03369_));
 sky130_fd_sc_hd__buf_8 _09030_ (.A(_03299_),
    .X(_03370_));
 sky130_fd_sc_hd__buf_6 _09031_ (.A(_02276_),
    .X(_03371_));
 sky130_fd_sc_hd__mux4_1 _09032_ (.A0(\regs[0][29] ),
    .A1(\regs[1][29] ),
    .A2(\regs[2][29] ),
    .A3(\regs[3][29] ),
    .S0(_03370_),
    .S1(_03371_),
    .X(_03372_));
 sky130_fd_sc_hd__mux4_1 _09033_ (.A0(\regs[4][29] ),
    .A1(\regs[5][29] ),
    .A2(\regs[6][29] ),
    .A3(\regs[7][29] ),
    .S0(_03370_),
    .S1(_03371_),
    .X(_03373_));
 sky130_fd_sc_hd__clkbuf_16 _09034_ (.A(_03243_),
    .X(_03374_));
 sky130_fd_sc_hd__mux2_1 _09035_ (.A0(_03372_),
    .A1(_03373_),
    .S(_03374_),
    .X(_03375_));
 sky130_fd_sc_hd__buf_6 _09036_ (.A(_03309_),
    .X(_03376_));
 sky130_fd_sc_hd__a221o_1 _09037_ (.A1(_03365_),
    .A2(_03369_),
    .B1(_03375_),
    .B2(_03376_),
    .C1(_03233_),
    .X(_03377_));
 sky130_fd_sc_hd__nor2_1 _09038_ (.A(_01693_),
    .B(_02993_),
    .Y(_03378_));
 sky130_fd_sc_hd__a31o_1 _09039_ (.A1(_00001_),
    .A2(_03361_),
    .A3(_03377_),
    .B1(_03378_),
    .X(_01341_));
 sky130_fd_sc_hd__mux2_1 _09040_ (.A0(\regs[30][28] ),
    .A1(\regs[31][28] ),
    .S(_03342_),
    .X(_03379_));
 sky130_fd_sc_hd__and2_1 _09041_ (.A(_03246_),
    .B(_03379_),
    .X(_03380_));
 sky130_fd_sc_hd__mux2_1 _09042_ (.A0(\regs[28][28] ),
    .A1(\regs[29][28] ),
    .S(_03342_),
    .X(_03381_));
 sky130_fd_sc_hd__a21o_1 _09043_ (.A1(_03282_),
    .A2(_03381_),
    .B1(_03235_),
    .X(_03382_));
 sky130_fd_sc_hd__or2b_1 _09044_ (.A(\regs[27][28] ),
    .B_N(_03280_),
    .X(_03383_));
 sky130_fd_sc_hd__buf_4 _09045_ (.A(_02280_),
    .X(_03384_));
 sky130_fd_sc_hd__o21a_1 _09046_ (.A1(_03384_),
    .A2(\regs[26][28] ),
    .B1(_03239_),
    .X(_03385_));
 sky130_fd_sc_hd__buf_6 _09047_ (.A(_02280_),
    .X(_03386_));
 sky130_fd_sc_hd__mux2_1 _09048_ (.A0(\regs[24][28] ),
    .A1(\regs[25][28] ),
    .S(_03386_),
    .X(_03387_));
 sky130_fd_sc_hd__a221o_1 _09049_ (.A1(_03383_),
    .A2(_03385_),
    .B1(_03387_),
    .B2(_03355_),
    .C1(_03254_),
    .X(_03388_));
 sky130_fd_sc_hd__o211a_1 _09050_ (.A1(_03380_),
    .A2(_03382_),
    .B1(_03388_),
    .C1(_03266_),
    .X(_03389_));
 sky130_fd_sc_hd__mux4_1 _09051_ (.A0(\regs[16][28] ),
    .A1(\regs[17][28] ),
    .A2(\regs[18][28] ),
    .A3(\regs[19][28] ),
    .S0(_03270_),
    .S1(_03304_),
    .X(_03390_));
 sky130_fd_sc_hd__mux4_1 _09052_ (.A0(\regs[20][28] ),
    .A1(\regs[21][28] ),
    .A2(\regs[22][28] ),
    .A3(\regs[23][28] ),
    .S0(_03269_),
    .S1(_03250_),
    .X(_03391_));
 sky130_fd_sc_hd__or2_1 _09053_ (.A(_03235_),
    .B(_03391_),
    .X(_03392_));
 sky130_fd_sc_hd__o211a_1 _09054_ (.A1(_02272_),
    .A2(_03390_),
    .B1(_03392_),
    .C1(_03258_),
    .X(_03393_));
 sky130_fd_sc_hd__buf_6 _09055_ (.A(_03235_),
    .X(_03394_));
 sky130_fd_sc_hd__buf_6 _09056_ (.A(_03245_),
    .X(_03395_));
 sky130_fd_sc_hd__mux4_1 _09057_ (.A0(\regs[12][28] ),
    .A1(\regs[13][28] ),
    .A2(\regs[14][28] ),
    .A3(\regs[15][28] ),
    .S0(_02282_),
    .S1(_03395_),
    .X(_03396_));
 sky130_fd_sc_hd__mux4_1 _09058_ (.A0(\regs[8][28] ),
    .A1(\regs[9][28] ),
    .A2(\regs[10][28] ),
    .A3(\regs[11][28] ),
    .S0(_02281_),
    .S1(_03245_),
    .X(_03397_));
 sky130_fd_sc_hd__or2_1 _09059_ (.A(_02271_),
    .B(_03397_),
    .X(_03398_));
 sky130_fd_sc_hd__o211a_1 _09060_ (.A1(_03394_),
    .A2(_03396_),
    .B1(_03398_),
    .C1(_03267_),
    .X(_03399_));
 sky130_fd_sc_hd__buf_8 _09061_ (.A(net14),
    .X(_03400_));
 sky130_fd_sc_hd__buf_6 _09062_ (.A(net15),
    .X(_03401_));
 sky130_fd_sc_hd__mux4_1 _09063_ (.A0(\regs[0][28] ),
    .A1(\regs[1][28] ),
    .A2(\regs[2][28] ),
    .A3(\regs[3][28] ),
    .S0(_03400_),
    .S1(_03401_),
    .X(_03402_));
 sky130_fd_sc_hd__mux4_1 _09064_ (.A0(\regs[4][28] ),
    .A1(\regs[5][28] ),
    .A2(\regs[6][28] ),
    .A3(\regs[7][28] ),
    .S0(_03237_),
    .S1(_03401_),
    .X(_03403_));
 sky130_fd_sc_hd__mux2_1 _09065_ (.A0(_03402_),
    .A1(_03403_),
    .S(_02271_),
    .X(_03404_));
 sky130_fd_sc_hd__a21o_1 _09066_ (.A1(_03309_),
    .A2(_03404_),
    .B1(_03233_),
    .X(_03405_));
 sky130_fd_sc_hd__o32a_1 _09067_ (.A1(_02264_),
    .A2(_03389_),
    .A3(_03393_),
    .B1(_03399_),
    .B2(_03405_),
    .X(_03406_));
 sky130_fd_sc_hd__mux2_1 _09068_ (.A0(\rs2_content[28] ),
    .A1(_03406_),
    .S(_02324_),
    .X(_03407_));
 sky130_fd_sc_hd__clkbuf_1 _09069_ (.A(_03407_),
    .X(_01340_));
 sky130_fd_sc_hd__buf_4 _09070_ (.A(_02255_),
    .X(_03408_));
 sky130_fd_sc_hd__mux4_1 _09071_ (.A0(\regs[12][27] ),
    .A1(\regs[13][27] ),
    .A2(\regs[14][27] ),
    .A3(\regs[15][27] ),
    .S0(_03290_),
    .S1(_03291_),
    .X(_03409_));
 sky130_fd_sc_hd__or2_1 _09072_ (.A(_03362_),
    .B(_03409_),
    .X(_03410_));
 sky130_fd_sc_hd__mux4_1 _09073_ (.A0(\regs[8][27] ),
    .A1(\regs[9][27] ),
    .A2(\regs[10][27] ),
    .A3(\regs[11][27] ),
    .S0(_03294_),
    .S1(_03295_),
    .X(_03411_));
 sky130_fd_sc_hd__o21a_1 _09074_ (.A1(_03316_),
    .A2(_03411_),
    .B1(_03297_),
    .X(_03412_));
 sky130_fd_sc_hd__mux4_1 _09075_ (.A0(\regs[0][27] ),
    .A1(\regs[1][27] ),
    .A2(\regs[2][27] ),
    .A3(\regs[3][27] ),
    .S0(_03300_),
    .S1(_03301_),
    .X(_03413_));
 sky130_fd_sc_hd__mux4_1 _09076_ (.A0(\regs[4][27] ),
    .A1(\regs[5][27] ),
    .A2(\regs[6][27] ),
    .A3(\regs[7][27] ),
    .S0(_03303_),
    .S1(_03305_),
    .X(_03414_));
 sky130_fd_sc_hd__mux2_1 _09077_ (.A0(_03413_),
    .A1(_03414_),
    .S(_03307_),
    .X(_03415_));
 sky130_fd_sc_hd__a22o_1 _09078_ (.A1(_03410_),
    .A2(_03412_),
    .B1(_03415_),
    .B2(_03310_),
    .X(_03416_));
 sky130_fd_sc_hd__mux4_1 _09079_ (.A0(\regs[16][27] ),
    .A1(\regs[17][27] ),
    .A2(\regs[18][27] ),
    .A3(\regs[19][27] ),
    .S0(_02283_),
    .S1(_03313_),
    .X(_03417_));
 sky130_fd_sc_hd__buf_8 _09080_ (.A(_03246_),
    .X(_03418_));
 sky130_fd_sc_hd__mux4_1 _09081_ (.A0(\regs[20][27] ),
    .A1(\regs[21][27] ),
    .A2(\regs[22][27] ),
    .A3(\regs[23][27] ),
    .S0(_02283_),
    .S1(_03418_),
    .X(_03419_));
 sky130_fd_sc_hd__mux2_1 _09082_ (.A0(_03417_),
    .A1(_03419_),
    .S(_03316_),
    .X(_03420_));
 sky130_fd_sc_hd__mux2_1 _09083_ (.A0(\regs[30][27] ),
    .A1(\regs[31][27] ),
    .S(_03318_),
    .X(_03421_));
 sky130_fd_sc_hd__mux2_1 _09084_ (.A0(\regs[28][27] ),
    .A1(\regs[29][27] ),
    .S(_03289_),
    .X(_03422_));
 sky130_fd_sc_hd__a21o_1 _09085_ (.A1(_03320_),
    .A2(_03422_),
    .B1(_03287_),
    .X(_03423_));
 sky130_fd_sc_hd__a21o_1 _09086_ (.A1(_02278_),
    .A2(_03421_),
    .B1(_03423_),
    .X(_03424_));
 sky130_fd_sc_hd__or2b_1 _09087_ (.A(\regs[27][27] ),
    .B_N(_03324_),
    .X(_03425_));
 sky130_fd_sc_hd__o21a_1 _09088_ (.A1(_03290_),
    .A2(\regs[26][27] ),
    .B1(_02277_),
    .X(_03426_));
 sky130_fd_sc_hd__mux2_1 _09089_ (.A0(\regs[24][27] ),
    .A1(\regs[25][27] ),
    .S(_03327_),
    .X(_03427_));
 sky130_fd_sc_hd__a221o_1 _09090_ (.A1(_03425_),
    .A2(_03426_),
    .B1(_03427_),
    .B2(_03329_),
    .C1(_03244_),
    .X(_03428_));
 sky130_fd_sc_hd__a31o_1 _09091_ (.A1(_02268_),
    .A2(_03424_),
    .A3(_03428_),
    .B1(_03331_),
    .X(_03429_));
 sky130_fd_sc_hd__a21o_1 _09092_ (.A1(_03312_),
    .A2(_03420_),
    .B1(_03429_),
    .X(_03430_));
 sky130_fd_sc_hd__o221a_1 _09093_ (.A1(\rs2_content[27] ),
    .A2(_03408_),
    .B1(_02266_),
    .B2(_03416_),
    .C1(_03430_),
    .X(_01339_));
 sky130_fd_sc_hd__mux4_1 _09094_ (.A0(\regs[16][26] ),
    .A1(\regs[17][26] ),
    .A2(\regs[18][26] ),
    .A3(\regs[19][26] ),
    .S0(_03335_),
    .S1(_03336_),
    .X(_03431_));
 sky130_fd_sc_hd__mux4_1 _09095_ (.A0(\regs[20][26] ),
    .A1(\regs[21][26] ),
    .A2(\regs[22][26] ),
    .A3(\regs[23][26] ),
    .S0(_03335_),
    .S1(_03336_),
    .X(_03432_));
 sky130_fd_sc_hd__mux2_1 _09096_ (.A0(_03431_),
    .A1(_03432_),
    .S(_03339_),
    .X(_03433_));
 sky130_fd_sc_hd__mux2_1 _09097_ (.A0(\regs[30][26] ),
    .A1(\regs[31][26] ),
    .S(_03343_),
    .X(_03434_));
 sky130_fd_sc_hd__and2_1 _09098_ (.A(_03341_),
    .B(_03434_),
    .X(_03435_));
 sky130_fd_sc_hd__mux2_1 _09099_ (.A0(\regs[28][26] ),
    .A1(\regs[29][26] ),
    .S(_03346_),
    .X(_03436_));
 sky130_fd_sc_hd__a21o_1 _09100_ (.A1(_03356_),
    .A2(_03436_),
    .B1(_03236_),
    .X(_03437_));
 sky130_fd_sc_hd__or2b_1 _09101_ (.A(\regs[27][26] ),
    .B_N(_03350_),
    .X(_03438_));
 sky130_fd_sc_hd__o21a_1 _09102_ (.A1(_03350_),
    .A2(\regs[26][26] ),
    .B1(_03352_),
    .X(_03439_));
 sky130_fd_sc_hd__mux2_1 _09103_ (.A0(\regs[24][26] ),
    .A1(\regs[25][26] ),
    .S(_03343_),
    .X(_03440_));
 sky130_fd_sc_hd__a221o_1 _09104_ (.A1(_03438_),
    .A2(_03439_),
    .B1(_03440_),
    .B2(_03356_),
    .C1(_03357_),
    .X(_03441_));
 sky130_fd_sc_hd__o211a_1 _09105_ (.A1(_03435_),
    .A2(_03437_),
    .B1(_03441_),
    .C1(_03359_),
    .X(_03442_));
 sky130_fd_sc_hd__a211o_1 _09106_ (.A1(_03334_),
    .A2(_03433_),
    .B1(_03442_),
    .C1(_02264_),
    .X(_03443_));
 sky130_fd_sc_hd__mux4_1 _09107_ (.A0(\regs[12][26] ),
    .A1(\regs[13][26] ),
    .A2(\regs[14][26] ),
    .A3(\regs[15][26] ),
    .S0(_03363_),
    .S1(_03268_),
    .X(_03444_));
 sky130_fd_sc_hd__or2_1 _09108_ (.A(_03362_),
    .B(_03444_),
    .X(_03445_));
 sky130_fd_sc_hd__mux4_1 _09109_ (.A0(\regs[8][26] ),
    .A1(\regs[9][26] ),
    .A2(\regs[10][26] ),
    .A3(\regs[11][26] ),
    .S0(_03300_),
    .S1(_03301_),
    .X(_03446_));
 sky130_fd_sc_hd__o21a_1 _09110_ (.A1(_03366_),
    .A2(_03446_),
    .B1(_03267_),
    .X(_03447_));
 sky130_fd_sc_hd__mux4_1 _09111_ (.A0(\regs[0][26] ),
    .A1(\regs[1][26] ),
    .A2(\regs[2][26] ),
    .A3(\regs[3][26] ),
    .S0(_03370_),
    .S1(_03371_),
    .X(_03448_));
 sky130_fd_sc_hd__mux4_1 _09112_ (.A0(\regs[4][26] ),
    .A1(\regs[5][26] ),
    .A2(\regs[6][26] ),
    .A3(\regs[7][26] ),
    .S0(_03370_),
    .S1(_03371_),
    .X(_03449_));
 sky130_fd_sc_hd__mux2_1 _09113_ (.A0(_03448_),
    .A1(_03449_),
    .S(_03374_),
    .X(_03450_));
 sky130_fd_sc_hd__a221o_1 _09114_ (.A1(_03445_),
    .A2(_03447_),
    .B1(_03450_),
    .B2(_03376_),
    .C1(_03233_),
    .X(_03451_));
 sky130_fd_sc_hd__nor2_1 _09115_ (.A(_01707_),
    .B(_02993_),
    .Y(_03452_));
 sky130_fd_sc_hd__a31o_1 _09116_ (.A1(_00001_),
    .A2(_03443_),
    .A3(_03451_),
    .B1(_03452_),
    .X(_01338_));
 sky130_fd_sc_hd__mux2_1 _09117_ (.A0(\regs[30][25] ),
    .A1(\regs[31][25] ),
    .S(_03386_),
    .X(_03453_));
 sky130_fd_sc_hd__and2_1 _09118_ (.A(_03246_),
    .B(_03453_),
    .X(_03454_));
 sky130_fd_sc_hd__mux2_1 _09119_ (.A0(\regs[28][25] ),
    .A1(\regs[29][25] ),
    .S(_03342_),
    .X(_03455_));
 sky130_fd_sc_hd__a21o_1 _09120_ (.A1(_03282_),
    .A2(_03455_),
    .B1(_03235_),
    .X(_03456_));
 sky130_fd_sc_hd__or2b_1 _09121_ (.A(\regs[27][25] ),
    .B_N(_03280_),
    .X(_03457_));
 sky130_fd_sc_hd__o21a_1 _09122_ (.A1(_03384_),
    .A2(\regs[26][25] ),
    .B1(_03239_),
    .X(_03458_));
 sky130_fd_sc_hd__mux2_1 _09123_ (.A0(\regs[24][25] ),
    .A1(\regs[25][25] ),
    .S(_03386_),
    .X(_03459_));
 sky130_fd_sc_hd__a221o_1 _09124_ (.A1(_03457_),
    .A2(_03458_),
    .B1(_03459_),
    .B2(_03355_),
    .C1(_03254_),
    .X(_03460_));
 sky130_fd_sc_hd__o211a_1 _09125_ (.A1(_03454_),
    .A2(_03456_),
    .B1(_03460_),
    .C1(_03266_),
    .X(_03461_));
 sky130_fd_sc_hd__mux4_1 _09126_ (.A0(\regs[16][25] ),
    .A1(\regs[17][25] ),
    .A2(\regs[18][25] ),
    .A3(\regs[19][25] ),
    .S0(_03270_),
    .S1(_03304_),
    .X(_03462_));
 sky130_fd_sc_hd__mux4_1 _09127_ (.A0(\regs[20][25] ),
    .A1(\regs[21][25] ),
    .A2(\regs[22][25] ),
    .A3(\regs[23][25] ),
    .S0(_03269_),
    .S1(_03250_),
    .X(_03463_));
 sky130_fd_sc_hd__or2_1 _09128_ (.A(_03274_),
    .B(_03463_),
    .X(_03464_));
 sky130_fd_sc_hd__o211a_1 _09129_ (.A1(_02272_),
    .A2(_03462_),
    .B1(_03464_),
    .C1(_03258_),
    .X(_03465_));
 sky130_fd_sc_hd__mux4_1 _09130_ (.A0(\regs[12][25] ),
    .A1(\regs[13][25] ),
    .A2(\regs[14][25] ),
    .A3(\regs[15][25] ),
    .S0(_02282_),
    .S1(_03395_),
    .X(_03466_));
 sky130_fd_sc_hd__mux4_1 _09131_ (.A0(\regs[8][25] ),
    .A1(\regs[9][25] ),
    .A2(\regs[10][25] ),
    .A3(\regs[11][25] ),
    .S0(_02281_),
    .S1(_03245_),
    .X(_03467_));
 sky130_fd_sc_hd__or2_1 _09132_ (.A(_02271_),
    .B(_03467_),
    .X(_03468_));
 sky130_fd_sc_hd__o211a_1 _09133_ (.A1(_03394_),
    .A2(_03466_),
    .B1(_03468_),
    .C1(_03267_),
    .X(_03469_));
 sky130_fd_sc_hd__mux4_1 _09134_ (.A0(\regs[0][25] ),
    .A1(\regs[1][25] ),
    .A2(\regs[2][25] ),
    .A3(\regs[3][25] ),
    .S0(_03400_),
    .S1(_03401_),
    .X(_03470_));
 sky130_fd_sc_hd__mux4_1 _09135_ (.A0(\regs[4][25] ),
    .A1(\regs[5][25] ),
    .A2(\regs[6][25] ),
    .A3(\regs[7][25] ),
    .S0(_03237_),
    .S1(_03401_),
    .X(_03471_));
 sky130_fd_sc_hd__mux2_1 _09136_ (.A0(_03470_),
    .A1(_03471_),
    .S(_03254_),
    .X(_03472_));
 sky130_fd_sc_hd__a21o_1 _09137_ (.A1(_03309_),
    .A2(_03472_),
    .B1(net18),
    .X(_03473_));
 sky130_fd_sc_hd__o32a_2 _09138_ (.A1(_02264_),
    .A2(_03461_),
    .A3(_03465_),
    .B1(_03469_),
    .B2(_03473_),
    .X(_03474_));
 sky130_fd_sc_hd__mux2_1 _09139_ (.A0(\rs2_content[25] ),
    .A1(_03474_),
    .S(_02253_),
    .X(_03475_));
 sky130_fd_sc_hd__clkbuf_1 _09140_ (.A(_03475_),
    .X(_01337_));
 sky130_fd_sc_hd__mux4_1 _09141_ (.A0(\regs[12][24] ),
    .A1(\regs[13][24] ),
    .A2(\regs[14][24] ),
    .A3(\regs[15][24] ),
    .S0(_03290_),
    .S1(_03291_),
    .X(_03476_));
 sky130_fd_sc_hd__or2_1 _09142_ (.A(_03362_),
    .B(_03476_),
    .X(_03477_));
 sky130_fd_sc_hd__mux4_1 _09143_ (.A0(\regs[8][24] ),
    .A1(\regs[9][24] ),
    .A2(\regs[10][24] ),
    .A3(\regs[11][24] ),
    .S0(_03294_),
    .S1(_03295_),
    .X(_03478_));
 sky130_fd_sc_hd__o21a_1 _09144_ (.A1(_03316_),
    .A2(_03478_),
    .B1(_03297_),
    .X(_03479_));
 sky130_fd_sc_hd__mux4_1 _09145_ (.A0(\regs[0][24] ),
    .A1(\regs[1][24] ),
    .A2(\regs[2][24] ),
    .A3(\regs[3][24] ),
    .S0(_03300_),
    .S1(_03301_),
    .X(_03480_));
 sky130_fd_sc_hd__mux4_1 _09146_ (.A0(\regs[4][24] ),
    .A1(\regs[5][24] ),
    .A2(\regs[6][24] ),
    .A3(\regs[7][24] ),
    .S0(_03303_),
    .S1(_03305_),
    .X(_03481_));
 sky130_fd_sc_hd__mux2_1 _09147_ (.A0(_03480_),
    .A1(_03481_),
    .S(_03307_),
    .X(_03482_));
 sky130_fd_sc_hd__a22o_1 _09148_ (.A1(_03477_),
    .A2(_03479_),
    .B1(_03482_),
    .B2(_03310_),
    .X(_03483_));
 sky130_fd_sc_hd__buf_8 _09149_ (.A(_03277_),
    .X(_03484_));
 sky130_fd_sc_hd__buf_6 _09150_ (.A(_03240_),
    .X(_03485_));
 sky130_fd_sc_hd__mux4_1 _09151_ (.A0(\regs[20][24] ),
    .A1(\regs[21][24] ),
    .A2(\regs[22][24] ),
    .A3(\regs[23][24] ),
    .S0(_03484_),
    .S1(_03485_),
    .X(_03486_));
 sky130_fd_sc_hd__buf_8 _09152_ (.A(_03277_),
    .X(_03487_));
 sky130_fd_sc_hd__buf_6 _09153_ (.A(_03240_),
    .X(_03488_));
 sky130_fd_sc_hd__mux4_1 _09154_ (.A0(\regs[16][24] ),
    .A1(\regs[17][24] ),
    .A2(\regs[18][24] ),
    .A3(\regs[19][24] ),
    .S0(_03487_),
    .S1(_03488_),
    .X(_03489_));
 sky130_fd_sc_hd__mux2_1 _09155_ (.A0(_03486_),
    .A1(_03489_),
    .S(_03394_),
    .X(_03490_));
 sky130_fd_sc_hd__mux2_1 _09156_ (.A0(\regs[30][24] ),
    .A1(\regs[31][24] ),
    .S(_03346_),
    .X(_03491_));
 sky130_fd_sc_hd__and2_1 _09157_ (.A(_03341_),
    .B(_03491_),
    .X(_03492_));
 sky130_fd_sc_hd__mux2_1 _09158_ (.A0(\regs[28][24] ),
    .A1(\regs[29][24] ),
    .S(_03327_),
    .X(_03493_));
 sky130_fd_sc_hd__a21o_1 _09159_ (.A1(_03329_),
    .A2(_03493_),
    .B1(_03394_),
    .X(_03494_));
 sky130_fd_sc_hd__or2b_1 _09160_ (.A(\regs[27][24] ),
    .B_N(_03363_),
    .X(_03495_));
 sky130_fd_sc_hd__o21a_1 _09161_ (.A1(_03363_),
    .A2(\regs[26][24] ),
    .B1(_03262_),
    .X(_03496_));
 sky130_fd_sc_hd__mux2_1 _09162_ (.A0(\regs[24][24] ),
    .A1(\regs[25][24] ),
    .S(_03346_),
    .X(_03497_));
 sky130_fd_sc_hd__a221o_1 _09163_ (.A1(_03495_),
    .A2(_03496_),
    .B1(_03497_),
    .B2(_03356_),
    .C1(_02272_),
    .X(_03498_));
 sky130_fd_sc_hd__o211a_1 _09164_ (.A1(_03492_),
    .A2(_03494_),
    .B1(_03498_),
    .C1(_02268_),
    .X(_03499_));
 sky130_fd_sc_hd__buf_6 _09165_ (.A(_03331_),
    .X(_03500_));
 sky130_fd_sc_hd__a211o_1 _09166_ (.A1(_03312_),
    .A2(_03490_),
    .B1(_03499_),
    .C1(_03500_),
    .X(_03501_));
 sky130_fd_sc_hd__o221a_1 _09167_ (.A1(\rs2_content[24] ),
    .A2(_03408_),
    .B1(_02266_),
    .B2(_03483_),
    .C1(_03501_),
    .X(_01336_));
 sky130_fd_sc_hd__mux2_1 _09168_ (.A0(\regs[30][23] ),
    .A1(\regs[31][23] ),
    .S(_03386_),
    .X(_03502_));
 sky130_fd_sc_hd__and2_1 _09169_ (.A(_03246_),
    .B(_03502_),
    .X(_03503_));
 sky130_fd_sc_hd__mux2_1 _09170_ (.A0(\regs[28][23] ),
    .A1(\regs[29][23] ),
    .S(_03342_),
    .X(_03504_));
 sky130_fd_sc_hd__a21o_1 _09171_ (.A1(_03282_),
    .A2(_03504_),
    .B1(_03235_),
    .X(_03505_));
 sky130_fd_sc_hd__or2b_1 _09172_ (.A(\regs[27][23] ),
    .B_N(_03280_),
    .X(_03506_));
 sky130_fd_sc_hd__o21a_1 _09173_ (.A1(_03384_),
    .A2(\regs[26][23] ),
    .B1(_03239_),
    .X(_03507_));
 sky130_fd_sc_hd__mux2_1 _09174_ (.A0(\regs[24][23] ),
    .A1(\regs[25][23] ),
    .S(_03386_),
    .X(_03508_));
 sky130_fd_sc_hd__a221o_1 _09175_ (.A1(_03506_),
    .A2(_03507_),
    .B1(_03508_),
    .B2(_03355_),
    .C1(_03254_),
    .X(_03509_));
 sky130_fd_sc_hd__o211a_1 _09176_ (.A1(_03503_),
    .A2(_03505_),
    .B1(_03509_),
    .C1(_03266_),
    .X(_03510_));
 sky130_fd_sc_hd__mux4_1 _09177_ (.A0(\regs[16][23] ),
    .A1(\regs[17][23] ),
    .A2(\regs[18][23] ),
    .A3(\regs[19][23] ),
    .S0(_03270_),
    .S1(_03304_),
    .X(_03511_));
 sky130_fd_sc_hd__mux4_1 _09178_ (.A0(\regs[20][23] ),
    .A1(\regs[21][23] ),
    .A2(\regs[22][23] ),
    .A3(\regs[23][23] ),
    .S0(_03269_),
    .S1(_03250_),
    .X(_03512_));
 sky130_fd_sc_hd__or2_1 _09179_ (.A(_03274_),
    .B(_03512_),
    .X(_03513_));
 sky130_fd_sc_hd__o211a_1 _09180_ (.A1(_03357_),
    .A2(_03511_),
    .B1(_03513_),
    .C1(_03258_),
    .X(_03514_));
 sky130_fd_sc_hd__mux4_1 _09181_ (.A0(\regs[12][23] ),
    .A1(\regs[13][23] ),
    .A2(\regs[14][23] ),
    .A3(\regs[15][23] ),
    .S0(_02282_),
    .S1(_03395_),
    .X(_03515_));
 sky130_fd_sc_hd__mux4_1 _09182_ (.A0(\regs[8][23] ),
    .A1(\regs[9][23] ),
    .A2(\regs[10][23] ),
    .A3(\regs[11][23] ),
    .S0(_02281_),
    .S1(_03245_),
    .X(_03516_));
 sky130_fd_sc_hd__or2_1 _09183_ (.A(_02271_),
    .B(_03516_),
    .X(_03517_));
 sky130_fd_sc_hd__o211a_1 _09184_ (.A1(_03236_),
    .A2(_03515_),
    .B1(_03517_),
    .C1(_03267_),
    .X(_03518_));
 sky130_fd_sc_hd__mux4_1 _09185_ (.A0(\regs[0][23] ),
    .A1(\regs[1][23] ),
    .A2(\regs[2][23] ),
    .A3(\regs[3][23] ),
    .S0(_03400_),
    .S1(_03401_),
    .X(_03519_));
 sky130_fd_sc_hd__mux4_1 _09186_ (.A0(\regs[4][23] ),
    .A1(\regs[5][23] ),
    .A2(\regs[6][23] ),
    .A3(\regs[7][23] ),
    .S0(_03237_),
    .S1(_03401_),
    .X(_03520_));
 sky130_fd_sc_hd__mux2_1 _09187_ (.A0(_03519_),
    .A1(_03520_),
    .S(_03254_),
    .X(_03521_));
 sky130_fd_sc_hd__a21o_1 _09188_ (.A1(_03309_),
    .A2(_03521_),
    .B1(net18),
    .X(_03522_));
 sky130_fd_sc_hd__o32a_2 _09189_ (.A1(_02264_),
    .A2(_03510_),
    .A3(_03514_),
    .B1(_03518_),
    .B2(_03522_),
    .X(_03523_));
 sky130_fd_sc_hd__mux2_1 _09190_ (.A0(\rs2_content[23] ),
    .A1(_03523_),
    .S(_02253_),
    .X(_03524_));
 sky130_fd_sc_hd__clkbuf_1 _09191_ (.A(_03524_),
    .X(_01335_));
 sky130_fd_sc_hd__mux4_1 _09192_ (.A0(\regs[12][22] ),
    .A1(\regs[13][22] ),
    .A2(\regs[14][22] ),
    .A3(\regs[15][22] ),
    .S0(_03290_),
    .S1(_03291_),
    .X(_03525_));
 sky130_fd_sc_hd__or2_1 _09193_ (.A(_03362_),
    .B(_03525_),
    .X(_03526_));
 sky130_fd_sc_hd__mux4_1 _09194_ (.A0(\regs[8][22] ),
    .A1(\regs[9][22] ),
    .A2(\regs[10][22] ),
    .A3(\regs[11][22] ),
    .S0(_03294_),
    .S1(_03295_),
    .X(_03527_));
 sky130_fd_sc_hd__o21a_1 _09195_ (.A1(_03316_),
    .A2(_03527_),
    .B1(_03297_),
    .X(_03528_));
 sky130_fd_sc_hd__mux4_1 _09196_ (.A0(\regs[0][22] ),
    .A1(\regs[1][22] ),
    .A2(\regs[2][22] ),
    .A3(\regs[3][22] ),
    .S0(_03303_),
    .S1(_03301_),
    .X(_03529_));
 sky130_fd_sc_hd__mux4_1 _09197_ (.A0(\regs[4][22] ),
    .A1(\regs[5][22] ),
    .A2(\regs[6][22] ),
    .A3(\regs[7][22] ),
    .S0(_03303_),
    .S1(_03305_),
    .X(_03530_));
 sky130_fd_sc_hd__mux2_1 _09198_ (.A0(_03529_),
    .A1(_03530_),
    .S(_03307_),
    .X(_03531_));
 sky130_fd_sc_hd__a22o_1 _09199_ (.A1(_03526_),
    .A2(_03528_),
    .B1(_03531_),
    .B2(_03310_),
    .X(_03532_));
 sky130_fd_sc_hd__mux4_1 _09200_ (.A0(\regs[16][22] ),
    .A1(\regs[17][22] ),
    .A2(\regs[18][22] ),
    .A3(\regs[19][22] ),
    .S0(_02283_),
    .S1(_03313_),
    .X(_03533_));
 sky130_fd_sc_hd__clkbuf_16 _09201_ (.A(_03238_),
    .X(_03534_));
 sky130_fd_sc_hd__mux4_1 _09202_ (.A0(\regs[20][22] ),
    .A1(\regs[21][22] ),
    .A2(\regs[22][22] ),
    .A3(\regs[23][22] ),
    .S0(_03534_),
    .S1(_03418_),
    .X(_03535_));
 sky130_fd_sc_hd__mux2_1 _09203_ (.A0(_03533_),
    .A1(_03535_),
    .S(_03366_),
    .X(_03536_));
 sky130_fd_sc_hd__or2b_1 _09204_ (.A(\regs[27][22] ),
    .B_N(_03324_),
    .X(_03537_));
 sky130_fd_sc_hd__o21a_1 _09205_ (.A1(_03324_),
    .A2(\regs[26][22] ),
    .B1(_02277_),
    .X(_03538_));
 sky130_fd_sc_hd__buf_4 _09206_ (.A(_03349_),
    .X(_03539_));
 sky130_fd_sc_hd__mux2_1 _09207_ (.A0(\regs[24][22] ),
    .A1(\regs[25][22] ),
    .S(_03539_),
    .X(_03540_));
 sky130_fd_sc_hd__a221o_1 _09208_ (.A1(_03537_),
    .A2(_03538_),
    .B1(_03540_),
    .B2(_03329_),
    .C1(_03374_),
    .X(_03541_));
 sky130_fd_sc_hd__mux2_1 _09209_ (.A0(\regs[30][22] ),
    .A1(\regs[31][22] ),
    .S(_03318_),
    .X(_03542_));
 sky130_fd_sc_hd__clkbuf_8 _09210_ (.A(_03272_),
    .X(_03543_));
 sky130_fd_sc_hd__mux2_1 _09211_ (.A0(\regs[28][22] ),
    .A1(\regs[29][22] ),
    .S(_03289_),
    .X(_03544_));
 sky130_fd_sc_hd__a21o_1 _09212_ (.A1(_03543_),
    .A2(_03544_),
    .B1(_03287_),
    .X(_03545_));
 sky130_fd_sc_hd__a21o_1 _09213_ (.A1(_02278_),
    .A2(_03542_),
    .B1(_03545_),
    .X(_03546_));
 sky130_fd_sc_hd__a31o_1 _09214_ (.A1(_02268_),
    .A2(_03541_),
    .A3(_03546_),
    .B1(_03331_),
    .X(_03547_));
 sky130_fd_sc_hd__a21o_1 _09215_ (.A1(_03312_),
    .A2(_03536_),
    .B1(_03547_),
    .X(_03548_));
 sky130_fd_sc_hd__o221a_1 _09216_ (.A1(\rs2_content[22] ),
    .A2(_03408_),
    .B1(_02266_),
    .B2(_03532_),
    .C1(_03548_),
    .X(_01334_));
 sky130_fd_sc_hd__mux4_1 _09217_ (.A0(\regs[0][21] ),
    .A1(\regs[1][21] ),
    .A2(\regs[2][21] ),
    .A3(\regs[3][21] ),
    .S0(_03363_),
    .S1(_03268_),
    .X(_03549_));
 sky130_fd_sc_hd__buf_8 _09218_ (.A(_03299_),
    .X(_03550_));
 sky130_fd_sc_hd__buf_8 _09219_ (.A(_02276_),
    .X(_03551_));
 sky130_fd_sc_hd__mux4_1 _09220_ (.A0(\regs[4][21] ),
    .A1(\regs[5][21] ),
    .A2(\regs[6][21] ),
    .A3(\regs[7][21] ),
    .S0(_03550_),
    .S1(_03551_),
    .X(_03552_));
 sky130_fd_sc_hd__mux2_1 _09221_ (.A0(_03549_),
    .A1(_03552_),
    .S(_03339_),
    .X(_03553_));
 sky130_fd_sc_hd__buf_8 _09222_ (.A(_03277_),
    .X(_03554_));
 sky130_fd_sc_hd__buf_6 _09223_ (.A(_03240_),
    .X(_03555_));
 sky130_fd_sc_hd__mux4_1 _09224_ (.A0(\regs[12][21] ),
    .A1(\regs[13][21] ),
    .A2(\regs[14][21] ),
    .A3(\regs[15][21] ),
    .S0(_03554_),
    .S1(_03555_),
    .X(_03556_));
 sky130_fd_sc_hd__or2_1 _09225_ (.A(_03288_),
    .B(_03556_),
    .X(_03557_));
 sky130_fd_sc_hd__mux4_1 _09226_ (.A0(\regs[8][21] ),
    .A1(\regs[9][21] ),
    .A2(\regs[10][21] ),
    .A3(\regs[11][21] ),
    .S0(_03534_),
    .S1(_03418_),
    .X(_03558_));
 sky130_fd_sc_hd__o21a_1 _09227_ (.A1(_02273_),
    .A2(_03558_),
    .B1(_03359_),
    .X(_03559_));
 sky130_fd_sc_hd__a22o_1 _09228_ (.A1(_03376_),
    .A2(_03553_),
    .B1(_03557_),
    .B2(_03559_),
    .X(_03560_));
 sky130_fd_sc_hd__mux4_1 _09229_ (.A0(\regs[16][21] ),
    .A1(\regs[17][21] ),
    .A2(\regs[18][21] ),
    .A3(\regs[19][21] ),
    .S0(_03484_),
    .S1(_03485_),
    .X(_03561_));
 sky130_fd_sc_hd__mux4_1 _09230_ (.A0(\regs[20][21] ),
    .A1(\regs[21][21] ),
    .A2(\regs[22][21] ),
    .A3(\regs[23][21] ),
    .S0(_03487_),
    .S1(_03488_),
    .X(_03562_));
 sky130_fd_sc_hd__mux2_1 _09231_ (.A0(_03561_),
    .A1(_03562_),
    .S(_03366_),
    .X(_03563_));
 sky130_fd_sc_hd__mux2_1 _09232_ (.A0(\regs[30][21] ),
    .A1(\regs[31][21] ),
    .S(_03327_),
    .X(_03564_));
 sky130_fd_sc_hd__mux2_1 _09233_ (.A0(\regs[28][21] ),
    .A1(\regs[29][21] ),
    .S(_03349_),
    .X(_03565_));
 sky130_fd_sc_hd__buf_6 _09234_ (.A(_03234_),
    .X(_03566_));
 sky130_fd_sc_hd__a21o_1 _09235_ (.A1(_03543_),
    .A2(_03565_),
    .B1(_03566_),
    .X(_03567_));
 sky130_fd_sc_hd__a21o_1 _09236_ (.A1(_02278_),
    .A2(_03564_),
    .B1(_03567_),
    .X(_03568_));
 sky130_fd_sc_hd__buf_4 _09237_ (.A(_03349_),
    .X(_03569_));
 sky130_fd_sc_hd__or2b_1 _09238_ (.A(\regs[27][21] ),
    .B_N(_03569_),
    .X(_03570_));
 sky130_fd_sc_hd__o21a_1 _09239_ (.A1(_03569_),
    .A2(\regs[26][21] ),
    .B1(_03352_),
    .X(_03571_));
 sky130_fd_sc_hd__mux2_1 _09240_ (.A0(\regs[24][21] ),
    .A1(\regs[25][21] ),
    .S(_03343_),
    .X(_03572_));
 sky130_fd_sc_hd__a221o_1 _09241_ (.A1(_03570_),
    .A2(_03571_),
    .B1(_03572_),
    .B2(_03356_),
    .C1(_03357_),
    .X(_03573_));
 sky130_fd_sc_hd__and3_1 _09242_ (.A(_03368_),
    .B(_03568_),
    .C(_03573_),
    .X(_03574_));
 sky130_fd_sc_hd__a211o_2 _09243_ (.A1(_03312_),
    .A2(_03563_),
    .B1(_03574_),
    .C1(_03500_),
    .X(_03575_));
 sky130_fd_sc_hd__o221a_1 _09244_ (.A1(\rs2_content[21] ),
    .A2(_03408_),
    .B1(_02266_),
    .B2(_03560_),
    .C1(_03575_),
    .X(_01333_));
 sky130_fd_sc_hd__mux4_1 _09245_ (.A0(\regs[12][20] ),
    .A1(\regs[13][20] ),
    .A2(\regs[14][20] ),
    .A3(\regs[15][20] ),
    .S0(_03238_),
    .S1(_03240_),
    .X(_03576_));
 sky130_fd_sc_hd__or2_1 _09246_ (.A(_03287_),
    .B(_03576_),
    .X(_03577_));
 sky130_fd_sc_hd__mux4_1 _09247_ (.A0(\regs[8][20] ),
    .A1(\regs[9][20] ),
    .A2(\regs[10][20] ),
    .A3(\regs[11][20] ),
    .S0(_03238_),
    .S1(_03246_),
    .X(_03578_));
 sky130_fd_sc_hd__o21a_1 _09248_ (.A1(_03244_),
    .A2(_03578_),
    .B1(_02267_),
    .X(_03579_));
 sky130_fd_sc_hd__mux4_1 _09249_ (.A0(\regs[0][20] ),
    .A1(\regs[1][20] ),
    .A2(\regs[2][20] ),
    .A3(\regs[3][20] ),
    .S0(_03249_),
    .S1(_03251_),
    .X(_03580_));
 sky130_fd_sc_hd__mux4_1 _09250_ (.A0(\regs[4][20] ),
    .A1(\regs[5][20] ),
    .A2(\regs[6][20] ),
    .A3(\regs[7][20] ),
    .S0(_03249_),
    .S1(_03251_),
    .X(_03581_));
 sky130_fd_sc_hd__mux2_1 _09251_ (.A0(_03580_),
    .A1(_03581_),
    .S(_03255_),
    .X(_03582_));
 sky130_fd_sc_hd__a22o_1 _09252_ (.A1(_03577_),
    .A2(_03579_),
    .B1(_03582_),
    .B2(_03259_),
    .X(_03583_));
 sky130_fd_sc_hd__mux4_1 _09253_ (.A0(\regs[16][20] ),
    .A1(\regs[17][20] ),
    .A2(\regs[18][20] ),
    .A3(\regs[19][20] ),
    .S0(_03261_),
    .S1(_03262_),
    .X(_03584_));
 sky130_fd_sc_hd__mux4_1 _09254_ (.A0(\regs[20][20] ),
    .A1(\regs[21][20] ),
    .A2(\regs[22][20] ),
    .A3(\regs[23][20] ),
    .S0(_02282_),
    .S1(_03262_),
    .X(_03585_));
 sky130_fd_sc_hd__mux2_1 _09255_ (.A0(_03584_),
    .A1(_03585_),
    .S(_02272_),
    .X(_03586_));
 sky130_fd_sc_hd__mux2_1 _09256_ (.A0(\regs[30][20] ),
    .A1(\regs[31][20] ),
    .S(_03270_),
    .X(_03587_));
 sky130_fd_sc_hd__mux2_1 _09257_ (.A0(\regs[28][20] ),
    .A1(\regs[29][20] ),
    .S(_03269_),
    .X(_03588_));
 sky130_fd_sc_hd__a21o_1 _09258_ (.A1(_03272_),
    .A2(_03588_),
    .B1(_03274_),
    .X(_03589_));
 sky130_fd_sc_hd__a21o_1 _09259_ (.A1(_03268_),
    .A2(_03587_),
    .B1(_03589_),
    .X(_03590_));
 sky130_fd_sc_hd__or2b_1 _09260_ (.A(\regs[27][20] ),
    .B_N(_03277_),
    .X(_03591_));
 sky130_fd_sc_hd__o21a_1 _09261_ (.A1(_03289_),
    .A2(\regs[26][20] ),
    .B1(_02276_),
    .X(_03592_));
 sky130_fd_sc_hd__mux2_1 _09262_ (.A0(\regs[24][20] ),
    .A1(\regs[25][20] ),
    .S(_03280_),
    .X(_03593_));
 sky130_fd_sc_hd__a221o_1 _09263_ (.A1(_03591_),
    .A2(_03592_),
    .B1(_03593_),
    .B2(_03282_),
    .C1(_03243_),
    .X(_03594_));
 sky130_fd_sc_hd__a31o_1 _09264_ (.A1(_03267_),
    .A2(_03590_),
    .A3(_03594_),
    .B1(_02263_),
    .X(_03595_));
 sky130_fd_sc_hd__a21o_1 _09265_ (.A1(_03259_),
    .A2(_03586_),
    .B1(_03595_),
    .X(_03596_));
 sky130_fd_sc_hd__o211a_2 _09266_ (.A1(_03233_),
    .A2(_03583_),
    .B1(_03596_),
    .C1(_02254_),
    .X(_03597_));
 sky130_fd_sc_hd__a21o_1 _09267_ (.A1(\rs2_content[20] ),
    .A2(_02543_),
    .B1(_03597_),
    .X(_01332_));
 sky130_fd_sc_hd__mux4_1 _09268_ (.A0(\regs[12][19] ),
    .A1(\regs[13][19] ),
    .A2(\regs[14][19] ),
    .A3(\regs[15][19] ),
    .S0(_03290_),
    .S1(_03291_),
    .X(_03598_));
 sky130_fd_sc_hd__or2_1 _09269_ (.A(_03362_),
    .B(_03598_),
    .X(_03599_));
 sky130_fd_sc_hd__mux4_1 _09270_ (.A0(\regs[8][19] ),
    .A1(\regs[9][19] ),
    .A2(\regs[10][19] ),
    .A3(\regs[11][19] ),
    .S0(_03294_),
    .S1(_03295_),
    .X(_03600_));
 sky130_fd_sc_hd__o21a_1 _09271_ (.A1(_03316_),
    .A2(_03600_),
    .B1(_03297_),
    .X(_03601_));
 sky130_fd_sc_hd__mux4_1 _09272_ (.A0(\regs[0][19] ),
    .A1(\regs[1][19] ),
    .A2(\regs[2][19] ),
    .A3(\regs[3][19] ),
    .S0(_03303_),
    .S1(_03301_),
    .X(_03602_));
 sky130_fd_sc_hd__mux4_1 _09273_ (.A0(\regs[4][19] ),
    .A1(\regs[5][19] ),
    .A2(\regs[6][19] ),
    .A3(\regs[7][19] ),
    .S0(_03318_),
    .S1(_03305_),
    .X(_03603_));
 sky130_fd_sc_hd__mux2_1 _09274_ (.A0(_03602_),
    .A1(_03603_),
    .S(_03339_),
    .X(_03604_));
 sky130_fd_sc_hd__a22o_1 _09275_ (.A1(_03599_),
    .A2(_03601_),
    .B1(_03604_),
    .B2(_03310_),
    .X(_03605_));
 sky130_fd_sc_hd__mux4_1 _09276_ (.A0(\regs[16][19] ),
    .A1(\regs[17][19] ),
    .A2(\regs[18][19] ),
    .A3(\regs[19][19] ),
    .S0(_02283_),
    .S1(_03313_),
    .X(_03606_));
 sky130_fd_sc_hd__mux4_1 _09277_ (.A0(\regs[20][19] ),
    .A1(\regs[21][19] ),
    .A2(\regs[22][19] ),
    .A3(\regs[23][19] ),
    .S0(_03534_),
    .S1(_03418_),
    .X(_03607_));
 sky130_fd_sc_hd__mux2_1 _09278_ (.A0(_03606_),
    .A1(_03607_),
    .S(_03366_),
    .X(_03608_));
 sky130_fd_sc_hd__or2b_1 _09279_ (.A(\regs[27][19] ),
    .B_N(_03324_),
    .X(_03609_));
 sky130_fd_sc_hd__o21a_1 _09280_ (.A1(_03324_),
    .A2(\regs[26][19] ),
    .B1(_02277_),
    .X(_03610_));
 sky130_fd_sc_hd__mux2_1 _09281_ (.A0(\regs[24][19] ),
    .A1(\regs[25][19] ),
    .S(_03539_),
    .X(_03611_));
 sky130_fd_sc_hd__a221o_1 _09282_ (.A1(_03609_),
    .A2(_03610_),
    .B1(_03611_),
    .B2(_03329_),
    .C1(_03244_),
    .X(_03612_));
 sky130_fd_sc_hd__mux2_1 _09283_ (.A0(\regs[30][19] ),
    .A1(\regs[31][19] ),
    .S(_03318_),
    .X(_03613_));
 sky130_fd_sc_hd__mux2_1 _09284_ (.A0(\regs[28][19] ),
    .A1(\regs[29][19] ),
    .S(_03289_),
    .X(_03614_));
 sky130_fd_sc_hd__a21o_1 _09285_ (.A1(_03543_),
    .A2(_03614_),
    .B1(_03287_),
    .X(_03615_));
 sky130_fd_sc_hd__a21o_1 _09286_ (.A1(_02278_),
    .A2(_03613_),
    .B1(_03615_),
    .X(_03616_));
 sky130_fd_sc_hd__a31o_1 _09287_ (.A1(_02268_),
    .A2(_03612_),
    .A3(_03616_),
    .B1(_03331_),
    .X(_03617_));
 sky130_fd_sc_hd__a21o_1 _09288_ (.A1(_03312_),
    .A2(_03608_),
    .B1(_03617_),
    .X(_03618_));
 sky130_fd_sc_hd__o221a_1 _09289_ (.A1(\rs2_content[19] ),
    .A2(_03408_),
    .B1(_02266_),
    .B2(_03605_),
    .C1(_03618_),
    .X(_01331_));
 sky130_fd_sc_hd__mux2_1 _09290_ (.A0(\regs[30][18] ),
    .A1(\regs[31][18] ),
    .S(_03386_),
    .X(_03619_));
 sky130_fd_sc_hd__and2_1 _09291_ (.A(_03246_),
    .B(_03619_),
    .X(_03620_));
 sky130_fd_sc_hd__mux2_1 _09292_ (.A0(\regs[28][18] ),
    .A1(\regs[29][18] ),
    .S(_03342_),
    .X(_03621_));
 sky130_fd_sc_hd__a21o_1 _09293_ (.A1(_03355_),
    .A2(_03621_),
    .B1(_03235_),
    .X(_03622_));
 sky130_fd_sc_hd__or2b_1 _09294_ (.A(\regs[27][18] ),
    .B_N(_03280_),
    .X(_03623_));
 sky130_fd_sc_hd__o21a_1 _09295_ (.A1(_03384_),
    .A2(\regs[26][18] ),
    .B1(_03239_),
    .X(_03624_));
 sky130_fd_sc_hd__mux2_1 _09296_ (.A0(\regs[24][18] ),
    .A1(\regs[25][18] ),
    .S(_02281_),
    .X(_03625_));
 sky130_fd_sc_hd__a221o_1 _09297_ (.A1(_03623_),
    .A2(_03624_),
    .B1(_03625_),
    .B2(_03355_),
    .C1(net16),
    .X(_03626_));
 sky130_fd_sc_hd__o211a_1 _09298_ (.A1(_03620_),
    .A2(_03622_),
    .B1(_03626_),
    .C1(_03266_),
    .X(_03627_));
 sky130_fd_sc_hd__mux4_1 _09299_ (.A0(\regs[16][18] ),
    .A1(\regs[17][18] ),
    .A2(\regs[18][18] ),
    .A3(\regs[19][18] ),
    .S0(_03270_),
    .S1(_03304_),
    .X(_03628_));
 sky130_fd_sc_hd__mux4_1 _09300_ (.A0(\regs[20][18] ),
    .A1(\regs[21][18] ),
    .A2(\regs[22][18] ),
    .A3(\regs[23][18] ),
    .S0(_03269_),
    .S1(_03250_),
    .X(_03629_));
 sky130_fd_sc_hd__or2_1 _09301_ (.A(_03274_),
    .B(_03629_),
    .X(_03630_));
 sky130_fd_sc_hd__o211a_1 _09302_ (.A1(_03357_),
    .A2(_03628_),
    .B1(_03630_),
    .C1(_03258_),
    .X(_03631_));
 sky130_fd_sc_hd__mux4_1 _09303_ (.A0(\regs[12][18] ),
    .A1(\regs[13][18] ),
    .A2(\regs[14][18] ),
    .A3(\regs[15][18] ),
    .S0(_02282_),
    .S1(_03395_),
    .X(_03632_));
 sky130_fd_sc_hd__mux4_1 _09304_ (.A0(\regs[8][18] ),
    .A1(\regs[9][18] ),
    .A2(\regs[10][18] ),
    .A3(\regs[11][18] ),
    .S0(_02281_),
    .S1(_03245_),
    .X(_03633_));
 sky130_fd_sc_hd__or2_1 _09305_ (.A(_02271_),
    .B(_03633_),
    .X(_03634_));
 sky130_fd_sc_hd__o211a_1 _09306_ (.A1(_03236_),
    .A2(_03632_),
    .B1(_03634_),
    .C1(_02267_),
    .X(_03635_));
 sky130_fd_sc_hd__mux4_1 _09307_ (.A0(\regs[0][18] ),
    .A1(\regs[1][18] ),
    .A2(\regs[2][18] ),
    .A3(\regs[3][18] ),
    .S0(_03400_),
    .S1(_03401_),
    .X(_03636_));
 sky130_fd_sc_hd__mux4_1 _09308_ (.A0(\regs[4][18] ),
    .A1(\regs[5][18] ),
    .A2(\regs[6][18] ),
    .A3(\regs[7][18] ),
    .S0(_03237_),
    .S1(_03239_),
    .X(_03637_));
 sky130_fd_sc_hd__mux2_1 _09309_ (.A0(_03636_),
    .A1(_03637_),
    .S(_03254_),
    .X(_03638_));
 sky130_fd_sc_hd__a21o_1 _09310_ (.A1(_03309_),
    .A2(_03638_),
    .B1(net18),
    .X(_03639_));
 sky130_fd_sc_hd__o32a_1 _09311_ (.A1(_02264_),
    .A2(_03627_),
    .A3(_03631_),
    .B1(_03635_),
    .B2(_03639_),
    .X(_03640_));
 sky130_fd_sc_hd__mux2_1 _09312_ (.A0(\rs2_content[18] ),
    .A1(_03640_),
    .S(_02253_),
    .X(_03641_));
 sky130_fd_sc_hd__clkbuf_1 _09313_ (.A(_03641_),
    .X(_01330_));
 sky130_fd_sc_hd__mux4_1 _09314_ (.A0(\regs[12][17] ),
    .A1(\regs[13][17] ),
    .A2(\regs[14][17] ),
    .A3(\regs[15][17] ),
    .S0(_03290_),
    .S1(_03291_),
    .X(_03642_));
 sky130_fd_sc_hd__or2_1 _09315_ (.A(_03362_),
    .B(_03642_),
    .X(_03643_));
 sky130_fd_sc_hd__mux4_2 _09316_ (.A0(\regs[8][17] ),
    .A1(\regs[9][17] ),
    .A2(\regs[10][17] ),
    .A3(\regs[11][17] ),
    .S0(_03294_),
    .S1(_03295_),
    .X(_03644_));
 sky130_fd_sc_hd__o21a_1 _09317_ (.A1(_03316_),
    .A2(_03644_),
    .B1(_03297_),
    .X(_03645_));
 sky130_fd_sc_hd__mux4_1 _09318_ (.A0(\regs[0][17] ),
    .A1(\regs[1][17] ),
    .A2(\regs[2][17] ),
    .A3(\regs[3][17] ),
    .S0(_03303_),
    .S1(_03301_),
    .X(_03646_));
 sky130_fd_sc_hd__mux4_1 _09319_ (.A0(\regs[4][17] ),
    .A1(\regs[5][17] ),
    .A2(\regs[6][17] ),
    .A3(\regs[7][17] ),
    .S0(_03318_),
    .S1(_03305_),
    .X(_03647_));
 sky130_fd_sc_hd__mux2_1 _09320_ (.A0(_03646_),
    .A1(_03647_),
    .S(_03339_),
    .X(_03648_));
 sky130_fd_sc_hd__a22o_1 _09321_ (.A1(_03643_),
    .A2(_03645_),
    .B1(_03648_),
    .B2(_03310_),
    .X(_03649_));
 sky130_fd_sc_hd__mux4_1 _09322_ (.A0(\regs[16][17] ),
    .A1(\regs[17][17] ),
    .A2(\regs[18][17] ),
    .A3(\regs[19][17] ),
    .S0(_02283_),
    .S1(_03313_),
    .X(_03650_));
 sky130_fd_sc_hd__mux4_1 _09323_ (.A0(\regs[20][17] ),
    .A1(\regs[21][17] ),
    .A2(\regs[22][17] ),
    .A3(\regs[23][17] ),
    .S0(_03534_),
    .S1(_03418_),
    .X(_03651_));
 sky130_fd_sc_hd__mux2_1 _09324_ (.A0(_03650_),
    .A1(_03651_),
    .S(_03366_),
    .X(_03652_));
 sky130_fd_sc_hd__or2b_1 _09325_ (.A(\regs[27][17] ),
    .B_N(_03324_),
    .X(_03653_));
 sky130_fd_sc_hd__o21a_1 _09326_ (.A1(_03324_),
    .A2(\regs[26][17] ),
    .B1(_02277_),
    .X(_03654_));
 sky130_fd_sc_hd__mux2_1 _09327_ (.A0(\regs[24][17] ),
    .A1(\regs[25][17] ),
    .S(_03539_),
    .X(_03655_));
 sky130_fd_sc_hd__a221o_1 _09328_ (.A1(_03653_),
    .A2(_03654_),
    .B1(_03655_),
    .B2(_03329_),
    .C1(_03244_),
    .X(_03656_));
 sky130_fd_sc_hd__mux2_1 _09329_ (.A0(\regs[30][17] ),
    .A1(\regs[31][17] ),
    .S(_03335_),
    .X(_03657_));
 sky130_fd_sc_hd__mux2_1 _09330_ (.A0(\regs[28][17] ),
    .A1(\regs[29][17] ),
    .S(_03289_),
    .X(_03658_));
 sky130_fd_sc_hd__a21o_1 _09331_ (.A1(_03543_),
    .A2(_03658_),
    .B1(_03566_),
    .X(_03659_));
 sky130_fd_sc_hd__a21o_1 _09332_ (.A1(_02278_),
    .A2(_03657_),
    .B1(_03659_),
    .X(_03660_));
 sky130_fd_sc_hd__a31o_1 _09333_ (.A1(_02268_),
    .A2(_03656_),
    .A3(_03660_),
    .B1(_03331_),
    .X(_03661_));
 sky130_fd_sc_hd__a21o_1 _09334_ (.A1(_03312_),
    .A2(_03652_),
    .B1(_03661_),
    .X(_03662_));
 sky130_fd_sc_hd__o221a_1 _09335_ (.A1(\rs2_content[17] ),
    .A2(_03408_),
    .B1(_02266_),
    .B2(_03649_),
    .C1(_03662_),
    .X(_01329_));
 sky130_fd_sc_hd__mux4_1 _09336_ (.A0(\regs[12][16] ),
    .A1(\regs[13][16] ),
    .A2(\regs[14][16] ),
    .A3(\regs[15][16] ),
    .S0(_03300_),
    .S1(_03291_),
    .X(_03663_));
 sky130_fd_sc_hd__or2_1 _09337_ (.A(_03362_),
    .B(_03663_),
    .X(_03664_));
 sky130_fd_sc_hd__mux4_1 _09338_ (.A0(\regs[8][16] ),
    .A1(\regs[9][16] ),
    .A2(\regs[10][16] ),
    .A3(\regs[11][16] ),
    .S0(_03294_),
    .S1(_03555_),
    .X(_03665_));
 sky130_fd_sc_hd__o21a_1 _09339_ (.A1(_03316_),
    .A2(_03665_),
    .B1(_03297_),
    .X(_03666_));
 sky130_fd_sc_hd__mux4_1 _09340_ (.A0(\regs[0][16] ),
    .A1(\regs[1][16] ),
    .A2(\regs[2][16] ),
    .A3(\regs[3][16] ),
    .S0(_03303_),
    .S1(_03305_),
    .X(_03667_));
 sky130_fd_sc_hd__mux4_1 _09341_ (.A0(\regs[4][16] ),
    .A1(\regs[5][16] ),
    .A2(\regs[6][16] ),
    .A3(\regs[7][16] ),
    .S0(_03318_),
    .S1(_03305_),
    .X(_03668_));
 sky130_fd_sc_hd__mux2_1 _09342_ (.A0(_03667_),
    .A1(_03668_),
    .S(_03339_),
    .X(_03669_));
 sky130_fd_sc_hd__a22o_1 _09343_ (.A1(_03664_),
    .A2(_03666_),
    .B1(_03669_),
    .B2(_03310_),
    .X(_03670_));
 sky130_fd_sc_hd__mux4_1 _09344_ (.A0(\regs[16][16] ),
    .A1(\regs[17][16] ),
    .A2(\regs[18][16] ),
    .A3(\regs[19][16] ),
    .S0(_02283_),
    .S1(_03313_),
    .X(_03671_));
 sky130_fd_sc_hd__mux4_1 _09345_ (.A0(\regs[20][16] ),
    .A1(\regs[21][16] ),
    .A2(\regs[22][16] ),
    .A3(\regs[23][16] ),
    .S0(_03534_),
    .S1(_03418_),
    .X(_03672_));
 sky130_fd_sc_hd__mux2_1 _09346_ (.A0(_03671_),
    .A1(_03672_),
    .S(_03366_),
    .X(_03673_));
 sky130_fd_sc_hd__mux2_1 _09347_ (.A0(\regs[30][16] ),
    .A1(\regs[31][16] ),
    .S(_03318_),
    .X(_03674_));
 sky130_fd_sc_hd__mux2_1 _09348_ (.A0(\regs[28][16] ),
    .A1(\regs[29][16] ),
    .S(_03289_),
    .X(_03675_));
 sky130_fd_sc_hd__a21o_1 _09349_ (.A1(_03320_),
    .A2(_03675_),
    .B1(_03287_),
    .X(_03676_));
 sky130_fd_sc_hd__a21o_1 _09350_ (.A1(_02278_),
    .A2(_03674_),
    .B1(_03676_),
    .X(_03677_));
 sky130_fd_sc_hd__or2b_1 _09351_ (.A(\regs[27][16] ),
    .B_N(_03290_),
    .X(_03678_));
 sky130_fd_sc_hd__o21a_1 _09352_ (.A1(_03290_),
    .A2(\regs[26][16] ),
    .B1(_02277_),
    .X(_03679_));
 sky130_fd_sc_hd__mux2_1 _09353_ (.A0(\regs[24][16] ),
    .A1(\regs[25][16] ),
    .S(_03327_),
    .X(_03680_));
 sky130_fd_sc_hd__a221o_1 _09354_ (.A1(_03678_),
    .A2(_03679_),
    .B1(_03680_),
    .B2(_03329_),
    .C1(_03244_),
    .X(_03681_));
 sky130_fd_sc_hd__a31o_1 _09355_ (.A1(_02268_),
    .A2(_03677_),
    .A3(_03681_),
    .B1(_03331_),
    .X(_03682_));
 sky130_fd_sc_hd__a21o_1 _09356_ (.A1(_03312_),
    .A2(_03673_),
    .B1(_03682_),
    .X(_03683_));
 sky130_fd_sc_hd__o221a_1 _09357_ (.A1(\rs2_content[16] ),
    .A2(_03408_),
    .B1(_02266_),
    .B2(_03670_),
    .C1(_03683_),
    .X(_01328_));
 sky130_fd_sc_hd__mux4_1 _09358_ (.A0(\regs[16][15] ),
    .A1(\regs[17][15] ),
    .A2(\regs[18][15] ),
    .A3(\regs[19][15] ),
    .S0(_03335_),
    .S1(_03336_),
    .X(_03684_));
 sky130_fd_sc_hd__mux4_1 _09359_ (.A0(\regs[20][15] ),
    .A1(\regs[21][15] ),
    .A2(\regs[22][15] ),
    .A3(\regs[23][15] ),
    .S0(_03335_),
    .S1(_03336_),
    .X(_03685_));
 sky130_fd_sc_hd__mux2_1 _09360_ (.A0(_03684_),
    .A1(_03685_),
    .S(_03339_),
    .X(_03686_));
 sky130_fd_sc_hd__mux2_1 _09361_ (.A0(\regs[30][15] ),
    .A1(\regs[31][15] ),
    .S(_03343_),
    .X(_03687_));
 sky130_fd_sc_hd__and2_1 _09362_ (.A(_03313_),
    .B(_03687_),
    .X(_03688_));
 sky130_fd_sc_hd__mux2_1 _09363_ (.A0(\regs[28][15] ),
    .A1(\regs[29][15] ),
    .S(_03346_),
    .X(_03689_));
 sky130_fd_sc_hd__a21o_1 _09364_ (.A1(_03356_),
    .A2(_03689_),
    .B1(_03236_),
    .X(_03690_));
 sky130_fd_sc_hd__or2b_1 _09365_ (.A(\regs[27][15] ),
    .B_N(_03350_),
    .X(_03691_));
 sky130_fd_sc_hd__o21a_1 _09366_ (.A1(_03350_),
    .A2(\regs[26][15] ),
    .B1(_03352_),
    .X(_03692_));
 sky130_fd_sc_hd__mux2_1 _09367_ (.A0(\regs[24][15] ),
    .A1(\regs[25][15] ),
    .S(_03343_),
    .X(_03693_));
 sky130_fd_sc_hd__a221o_1 _09368_ (.A1(_03691_),
    .A2(_03692_),
    .B1(_03693_),
    .B2(_03356_),
    .C1(_03357_),
    .X(_03694_));
 sky130_fd_sc_hd__o211a_1 _09369_ (.A1(_03688_),
    .A2(_03690_),
    .B1(_03694_),
    .C1(_03297_),
    .X(_03695_));
 sky130_fd_sc_hd__a211o_1 _09370_ (.A1(_03334_),
    .A2(_03686_),
    .B1(_03695_),
    .C1(_02264_),
    .X(_03696_));
 sky130_fd_sc_hd__mux4_1 _09371_ (.A0(\regs[12][15] ),
    .A1(\regs[13][15] ),
    .A2(\regs[14][15] ),
    .A3(\regs[15][15] ),
    .S0(_03363_),
    .S1(_03268_),
    .X(_03697_));
 sky130_fd_sc_hd__or2_1 _09372_ (.A(_03394_),
    .B(_03697_),
    .X(_03698_));
 sky130_fd_sc_hd__mux4_1 _09373_ (.A0(\regs[8][15] ),
    .A1(\regs[9][15] ),
    .A2(\regs[10][15] ),
    .A3(\regs[11][15] ),
    .S0(_03300_),
    .S1(_03301_),
    .X(_03699_));
 sky130_fd_sc_hd__o21a_1 _09374_ (.A1(_03366_),
    .A2(_03699_),
    .B1(_03267_),
    .X(_03700_));
 sky130_fd_sc_hd__mux4_1 _09375_ (.A0(\regs[0][15] ),
    .A1(\regs[1][15] ),
    .A2(\regs[2][15] ),
    .A3(\regs[3][15] ),
    .S0(_03370_),
    .S1(_03371_),
    .X(_03701_));
 sky130_fd_sc_hd__mux4_1 _09376_ (.A0(\regs[4][15] ),
    .A1(\regs[5][15] ),
    .A2(\regs[6][15] ),
    .A3(\regs[7][15] ),
    .S0(_03350_),
    .S1(_02277_),
    .X(_03702_));
 sky130_fd_sc_hd__mux2_1 _09377_ (.A0(_03701_),
    .A1(_03702_),
    .S(_03374_),
    .X(_03703_));
 sky130_fd_sc_hd__a221o_1 _09378_ (.A1(_03698_),
    .A2(_03700_),
    .B1(_03703_),
    .B2(_03259_),
    .C1(_03233_),
    .X(_03704_));
 sky130_fd_sc_hd__nor2_1 _09379_ (.A(_01741_),
    .B(_02993_),
    .Y(_03705_));
 sky130_fd_sc_hd__a31o_1 _09380_ (.A1(_00001_),
    .A2(_03696_),
    .A3(_03704_),
    .B1(_03705_),
    .X(_01327_));
 sky130_fd_sc_hd__mux4_1 _09381_ (.A0(\regs[0][14] ),
    .A1(\regs[1][14] ),
    .A2(\regs[2][14] ),
    .A3(\regs[3][14] ),
    .S0(_03363_),
    .S1(_03268_),
    .X(_03706_));
 sky130_fd_sc_hd__mux4_1 _09382_ (.A0(\regs[4][14] ),
    .A1(\regs[5][14] ),
    .A2(\regs[6][14] ),
    .A3(\regs[7][14] ),
    .S0(_03550_),
    .S1(_03551_),
    .X(_03707_));
 sky130_fd_sc_hd__mux2_1 _09383_ (.A0(_03706_),
    .A1(_03707_),
    .S(_03374_),
    .X(_03708_));
 sky130_fd_sc_hd__mux4_1 _09384_ (.A0(\regs[12][14] ),
    .A1(\regs[13][14] ),
    .A2(\regs[14][14] ),
    .A3(\regs[15][14] ),
    .S0(_03554_),
    .S1(_03555_),
    .X(_03709_));
 sky130_fd_sc_hd__or2_1 _09385_ (.A(_03288_),
    .B(_03709_),
    .X(_03710_));
 sky130_fd_sc_hd__mux4_1 _09386_ (.A0(\regs[8][14] ),
    .A1(\regs[9][14] ),
    .A2(\regs[10][14] ),
    .A3(\regs[11][14] ),
    .S0(_03534_),
    .S1(_03418_),
    .X(_03711_));
 sky130_fd_sc_hd__o21a_1 _09387_ (.A1(_02273_),
    .A2(_03711_),
    .B1(_03359_),
    .X(_03712_));
 sky130_fd_sc_hd__a22o_1 _09388_ (.A1(_03376_),
    .A2(_03708_),
    .B1(_03710_),
    .B2(_03712_),
    .X(_03713_));
 sky130_fd_sc_hd__mux4_1 _09389_ (.A0(\regs[16][14] ),
    .A1(\regs[17][14] ),
    .A2(\regs[18][14] ),
    .A3(\regs[19][14] ),
    .S0(_03484_),
    .S1(_03485_),
    .X(_03714_));
 sky130_fd_sc_hd__mux4_1 _09390_ (.A0(\regs[20][14] ),
    .A1(\regs[21][14] ),
    .A2(\regs[22][14] ),
    .A3(\regs[23][14] ),
    .S0(_03487_),
    .S1(_03488_),
    .X(_03715_));
 sky130_fd_sc_hd__mux2_1 _09391_ (.A0(_03714_),
    .A1(_03715_),
    .S(_03366_),
    .X(_03716_));
 sky130_fd_sc_hd__mux2_1 _09392_ (.A0(\regs[30][14] ),
    .A1(\regs[31][14] ),
    .S(_03327_),
    .X(_03717_));
 sky130_fd_sc_hd__mux2_1 _09393_ (.A0(\regs[28][14] ),
    .A1(\regs[29][14] ),
    .S(_03349_),
    .X(_03718_));
 sky130_fd_sc_hd__a21o_1 _09394_ (.A1(_03543_),
    .A2(_03718_),
    .B1(_03566_),
    .X(_03719_));
 sky130_fd_sc_hd__a21o_1 _09395_ (.A1(_02278_),
    .A2(_03717_),
    .B1(_03719_),
    .X(_03720_));
 sky130_fd_sc_hd__or2b_1 _09396_ (.A(\regs[27][14] ),
    .B_N(_03569_),
    .X(_03721_));
 sky130_fd_sc_hd__o21a_1 _09397_ (.A1(_03569_),
    .A2(\regs[26][14] ),
    .B1(_03352_),
    .X(_03722_));
 sky130_fd_sc_hd__mux2_1 _09398_ (.A0(\regs[24][14] ),
    .A1(\regs[25][14] ),
    .S(_03261_),
    .X(_03723_));
 sky130_fd_sc_hd__a221o_1 _09399_ (.A1(_03721_),
    .A2(_03722_),
    .B1(_03723_),
    .B2(_03320_),
    .C1(_03255_),
    .X(_03724_));
 sky130_fd_sc_hd__and3_1 _09400_ (.A(_03368_),
    .B(_03720_),
    .C(_03724_),
    .X(_03725_));
 sky130_fd_sc_hd__a211o_1 _09401_ (.A1(_03312_),
    .A2(_03716_),
    .B1(_03725_),
    .C1(_03500_),
    .X(_03726_));
 sky130_fd_sc_hd__o221a_1 _09402_ (.A1(\rs2_content[14] ),
    .A2(_03408_),
    .B1(_02266_),
    .B2(_03713_),
    .C1(_03726_),
    .X(_01326_));
 sky130_fd_sc_hd__mux4_1 _09403_ (.A0(\regs[12][13] ),
    .A1(\regs[13][13] ),
    .A2(\regs[14][13] ),
    .A3(\regs[15][13] ),
    .S0(_03249_),
    .S1(_03240_),
    .X(_03727_));
 sky130_fd_sc_hd__or2_1 _09404_ (.A(_03287_),
    .B(_03727_),
    .X(_03728_));
 sky130_fd_sc_hd__mux4_1 _09405_ (.A0(\regs[8][13] ),
    .A1(\regs[9][13] ),
    .A2(\regs[10][13] ),
    .A3(\regs[11][13] ),
    .S0(_03238_),
    .S1(_03246_),
    .X(_03729_));
 sky130_fd_sc_hd__o21a_1 _09406_ (.A1(_03244_),
    .A2(_03729_),
    .B1(_02267_),
    .X(_03730_));
 sky130_fd_sc_hd__mux4_1 _09407_ (.A0(\regs[0][13] ),
    .A1(\regs[1][13] ),
    .A2(\regs[2][13] ),
    .A3(\regs[3][13] ),
    .S0(_03249_),
    .S1(_03251_),
    .X(_03731_));
 sky130_fd_sc_hd__mux4_1 _09408_ (.A0(\regs[4][13] ),
    .A1(\regs[5][13] ),
    .A2(\regs[6][13] ),
    .A3(\regs[7][13] ),
    .S0(_03249_),
    .S1(_03251_),
    .X(_03732_));
 sky130_fd_sc_hd__mux2_1 _09409_ (.A0(_03731_),
    .A1(_03732_),
    .S(_03243_),
    .X(_03733_));
 sky130_fd_sc_hd__a22o_1 _09410_ (.A1(_03728_),
    .A2(_03730_),
    .B1(_03733_),
    .B2(_03259_),
    .X(_03734_));
 sky130_fd_sc_hd__mux4_1 _09411_ (.A0(\regs[16][13] ),
    .A1(\regs[17][13] ),
    .A2(\regs[18][13] ),
    .A3(\regs[19][13] ),
    .S0(_03261_),
    .S1(_03262_),
    .X(_03735_));
 sky130_fd_sc_hd__mux4_1 _09412_ (.A0(\regs[20][13] ),
    .A1(\regs[21][13] ),
    .A2(\regs[22][13] ),
    .A3(\regs[23][13] ),
    .S0(_02282_),
    .S1(_03262_),
    .X(_03736_));
 sky130_fd_sc_hd__mux2_1 _09413_ (.A0(_03735_),
    .A1(_03736_),
    .S(_02272_),
    .X(_03737_));
 sky130_fd_sc_hd__mux2_1 _09414_ (.A0(\regs[30][13] ),
    .A1(\regs[31][13] ),
    .S(_03299_),
    .X(_03738_));
 sky130_fd_sc_hd__mux2_1 _09415_ (.A0(\regs[28][13] ),
    .A1(\regs[29][13] ),
    .S(_03269_),
    .X(_03739_));
 sky130_fd_sc_hd__a21o_1 _09416_ (.A1(_03272_),
    .A2(_03739_),
    .B1(_03274_),
    .X(_03740_));
 sky130_fd_sc_hd__a21o_1 _09417_ (.A1(_03268_),
    .A2(_03738_),
    .B1(_03740_),
    .X(_03741_));
 sky130_fd_sc_hd__or2b_1 _09418_ (.A(\regs[27][13] ),
    .B_N(_03277_),
    .X(_03742_));
 sky130_fd_sc_hd__o21a_1 _09419_ (.A1(_03289_),
    .A2(\regs[26][13] ),
    .B1(_02276_),
    .X(_03743_));
 sky130_fd_sc_hd__mux2_1 _09420_ (.A0(\regs[24][13] ),
    .A1(\regs[25][13] ),
    .S(_03280_),
    .X(_03744_));
 sky130_fd_sc_hd__a221o_1 _09421_ (.A1(_03742_),
    .A2(_03743_),
    .B1(_03744_),
    .B2(_03282_),
    .C1(_03243_),
    .X(_03745_));
 sky130_fd_sc_hd__a31o_1 _09422_ (.A1(_03267_),
    .A2(_03741_),
    .A3(_03745_),
    .B1(_02263_),
    .X(_03746_));
 sky130_fd_sc_hd__a21o_1 _09423_ (.A1(_03259_),
    .A2(_03737_),
    .B1(_03746_),
    .X(_03747_));
 sky130_fd_sc_hd__o211a_1 _09424_ (.A1(_03233_),
    .A2(_03734_),
    .B1(_03747_),
    .C1(_02254_),
    .X(_03748_));
 sky130_fd_sc_hd__a21o_1 _09425_ (.A1(\rs2_content[13] ),
    .A2(_02543_),
    .B1(_03748_),
    .X(_01325_));
 sky130_fd_sc_hd__mux4_1 _09426_ (.A0(\regs[0][12] ),
    .A1(\regs[1][12] ),
    .A2(\regs[2][12] ),
    .A3(\regs[3][12] ),
    .S0(_03550_),
    .S1(_03551_),
    .X(_03749_));
 sky130_fd_sc_hd__mux4_1 _09427_ (.A0(\regs[4][12] ),
    .A1(\regs[5][12] ),
    .A2(\regs[6][12] ),
    .A3(\regs[7][12] ),
    .S0(_03550_),
    .S1(_03551_),
    .X(_03750_));
 sky130_fd_sc_hd__mux2_1 _09428_ (.A0(_03749_),
    .A1(_03750_),
    .S(_03374_),
    .X(_03751_));
 sky130_fd_sc_hd__mux4_1 _09429_ (.A0(\regs[12][12] ),
    .A1(\regs[13][12] ),
    .A2(\regs[14][12] ),
    .A3(\regs[15][12] ),
    .S0(_03554_),
    .S1(_03555_),
    .X(_03752_));
 sky130_fd_sc_hd__or2_1 _09430_ (.A(_03288_),
    .B(_03752_),
    .X(_03753_));
 sky130_fd_sc_hd__mux4_1 _09431_ (.A0(\regs[8][12] ),
    .A1(\regs[9][12] ),
    .A2(\regs[10][12] ),
    .A3(\regs[11][12] ),
    .S0(_03534_),
    .S1(_03418_),
    .X(_03754_));
 sky130_fd_sc_hd__o21a_1 _09432_ (.A1(_02273_),
    .A2(_03754_),
    .B1(_03359_),
    .X(_03755_));
 sky130_fd_sc_hd__a22o_1 _09433_ (.A1(_03376_),
    .A2(_03751_),
    .B1(_03753_),
    .B2(_03755_),
    .X(_03756_));
 sky130_fd_sc_hd__mux4_1 _09434_ (.A0(\regs[16][12] ),
    .A1(\regs[17][12] ),
    .A2(\regs[18][12] ),
    .A3(\regs[19][12] ),
    .S0(_03484_),
    .S1(_03485_),
    .X(_03757_));
 sky130_fd_sc_hd__mux4_1 _09435_ (.A0(\regs[20][12] ),
    .A1(\regs[21][12] ),
    .A2(\regs[22][12] ),
    .A3(\regs[23][12] ),
    .S0(_03487_),
    .S1(_03488_),
    .X(_03758_));
 sky130_fd_sc_hd__mux2_1 _09436_ (.A0(_03757_),
    .A1(_03758_),
    .S(_03307_),
    .X(_03759_));
 sky130_fd_sc_hd__mux2_1 _09437_ (.A0(\regs[30][12] ),
    .A1(\regs[31][12] ),
    .S(_03327_),
    .X(_03760_));
 sky130_fd_sc_hd__mux2_1 _09438_ (.A0(\regs[28][12] ),
    .A1(\regs[29][12] ),
    .S(_03349_),
    .X(_03761_));
 sky130_fd_sc_hd__a21o_1 _09439_ (.A1(_03543_),
    .A2(_03761_),
    .B1(_03566_),
    .X(_03762_));
 sky130_fd_sc_hd__a21o_1 _09440_ (.A1(_03341_),
    .A2(_03760_),
    .B1(_03762_),
    .X(_03763_));
 sky130_fd_sc_hd__or2b_1 _09441_ (.A(\regs[27][12] ),
    .B_N(_03569_),
    .X(_03764_));
 sky130_fd_sc_hd__o21a_1 _09442_ (.A1(_03539_),
    .A2(\regs[26][12] ),
    .B1(_03352_),
    .X(_03765_));
 sky130_fd_sc_hd__mux2_1 _09443_ (.A0(\regs[24][12] ),
    .A1(\regs[25][12] ),
    .S(_03261_),
    .X(_03766_));
 sky130_fd_sc_hd__a221o_1 _09444_ (.A1(_03764_),
    .A2(_03765_),
    .B1(_03766_),
    .B2(_03320_),
    .C1(_03255_),
    .X(_03767_));
 sky130_fd_sc_hd__and3_1 _09445_ (.A(_03368_),
    .B(_03763_),
    .C(_03767_),
    .X(_03768_));
 sky130_fd_sc_hd__a211o_1 _09446_ (.A1(_03334_),
    .A2(_03759_),
    .B1(_03768_),
    .C1(_03500_),
    .X(_03769_));
 sky130_fd_sc_hd__o221a_1 _09447_ (.A1(\rs2_content[12] ),
    .A2(_03408_),
    .B1(_02265_),
    .B2(_03756_),
    .C1(_03769_),
    .X(_01324_));
 sky130_fd_sc_hd__mux4_1 _09448_ (.A0(\regs[4][11] ),
    .A1(\regs[5][11] ),
    .A2(\regs[6][11] ),
    .A3(\regs[7][11] ),
    .S0(_03550_),
    .S1(_03551_),
    .X(_03770_));
 sky130_fd_sc_hd__mux4_1 _09449_ (.A0(\regs[0][11] ),
    .A1(\regs[1][11] ),
    .A2(\regs[2][11] ),
    .A3(\regs[3][11] ),
    .S0(_03550_),
    .S1(_03551_),
    .X(_03771_));
 sky130_fd_sc_hd__mux2_1 _09450_ (.A0(_03770_),
    .A1(_03771_),
    .S(_03394_),
    .X(_03772_));
 sky130_fd_sc_hd__mux4_1 _09451_ (.A0(\regs[12][11] ),
    .A1(\regs[13][11] ),
    .A2(\regs[14][11] ),
    .A3(\regs[15][11] ),
    .S0(_03554_),
    .S1(_03555_),
    .X(_03773_));
 sky130_fd_sc_hd__or2_1 _09452_ (.A(_03288_),
    .B(_03773_),
    .X(_03774_));
 sky130_fd_sc_hd__mux4_1 _09453_ (.A0(\regs[8][11] ),
    .A1(\regs[9][11] ),
    .A2(\regs[10][11] ),
    .A3(\regs[11][11] ),
    .S0(_03534_),
    .S1(_03418_),
    .X(_03775_));
 sky130_fd_sc_hd__o21a_1 _09454_ (.A1(_02273_),
    .A2(_03775_),
    .B1(_03359_),
    .X(_03776_));
 sky130_fd_sc_hd__a22o_1 _09455_ (.A1(_03376_),
    .A2(_03772_),
    .B1(_03774_),
    .B2(_03776_),
    .X(_03777_));
 sky130_fd_sc_hd__mux4_1 _09456_ (.A0(\regs[16][11] ),
    .A1(\regs[17][11] ),
    .A2(\regs[18][11] ),
    .A3(\regs[19][11] ),
    .S0(_03484_),
    .S1(_03485_),
    .X(_03778_));
 sky130_fd_sc_hd__mux4_1 _09457_ (.A0(\regs[20][11] ),
    .A1(\regs[21][11] ),
    .A2(\regs[22][11] ),
    .A3(\regs[23][11] ),
    .S0(_03487_),
    .S1(_03488_),
    .X(_03779_));
 sky130_fd_sc_hd__mux2_1 _09458_ (.A0(_03778_),
    .A1(_03779_),
    .S(_03307_),
    .X(_03780_));
 sky130_fd_sc_hd__mux2_1 _09459_ (.A0(\regs[30][11] ),
    .A1(\regs[31][11] ),
    .S(_03327_),
    .X(_03781_));
 sky130_fd_sc_hd__mux2_1 _09460_ (.A0(\regs[28][11] ),
    .A1(\regs[29][11] ),
    .S(_03349_),
    .X(_03782_));
 sky130_fd_sc_hd__a21o_1 _09461_ (.A1(_03543_),
    .A2(_03782_),
    .B1(_03566_),
    .X(_03783_));
 sky130_fd_sc_hd__a21o_1 _09462_ (.A1(_03341_),
    .A2(_03781_),
    .B1(_03783_),
    .X(_03784_));
 sky130_fd_sc_hd__or2b_1 _09463_ (.A(\regs[27][11] ),
    .B_N(_03569_),
    .X(_03785_));
 sky130_fd_sc_hd__o21a_1 _09464_ (.A1(_03539_),
    .A2(\regs[26][11] ),
    .B1(_03352_),
    .X(_03786_));
 sky130_fd_sc_hd__mux2_1 _09465_ (.A0(\regs[24][11] ),
    .A1(\regs[25][11] ),
    .S(_03261_),
    .X(_03787_));
 sky130_fd_sc_hd__a221o_1 _09466_ (.A1(_03785_),
    .A2(_03786_),
    .B1(_03787_),
    .B2(_03320_),
    .C1(_03255_),
    .X(_03788_));
 sky130_fd_sc_hd__and3_1 _09467_ (.A(_03368_),
    .B(_03784_),
    .C(_03788_),
    .X(_03789_));
 sky130_fd_sc_hd__a211o_1 _09468_ (.A1(_03334_),
    .A2(_03780_),
    .B1(_03789_),
    .C1(_03500_),
    .X(_03790_));
 sky130_fd_sc_hd__o221a_1 _09469_ (.A1(\rs2_content[11] ),
    .A2(_03408_),
    .B1(_02265_),
    .B2(_03777_),
    .C1(_03790_),
    .X(_01323_));
 sky130_fd_sc_hd__mux2_1 _09470_ (.A0(\regs[30][10] ),
    .A1(\regs[31][10] ),
    .S(_03386_),
    .X(_03791_));
 sky130_fd_sc_hd__and2_1 _09471_ (.A(_03246_),
    .B(_03791_),
    .X(_03792_));
 sky130_fd_sc_hd__mux2_1 _09472_ (.A0(\regs[28][10] ),
    .A1(\regs[29][10] ),
    .S(_03342_),
    .X(_03793_));
 sky130_fd_sc_hd__a21o_1 _09473_ (.A1(_03355_),
    .A2(_03793_),
    .B1(_03235_),
    .X(_03794_));
 sky130_fd_sc_hd__or2b_1 _09474_ (.A(\regs[27][10] ),
    .B_N(_03384_),
    .X(_03795_));
 sky130_fd_sc_hd__o21a_1 _09475_ (.A1(_03384_),
    .A2(\regs[26][10] ),
    .B1(_03250_),
    .X(_03796_));
 sky130_fd_sc_hd__mux2_1 _09476_ (.A0(\regs[24][10] ),
    .A1(\regs[25][10] ),
    .S(_02281_),
    .X(_03797_));
 sky130_fd_sc_hd__a221o_1 _09477_ (.A1(_03795_),
    .A2(_03796_),
    .B1(_03797_),
    .B2(_03355_),
    .C1(net16),
    .X(_03798_));
 sky130_fd_sc_hd__o211a_1 _09478_ (.A1(_03792_),
    .A2(_03794_),
    .B1(_03798_),
    .C1(_03266_),
    .X(_03799_));
 sky130_fd_sc_hd__mux4_1 _09479_ (.A0(\regs[16][10] ),
    .A1(\regs[17][10] ),
    .A2(\regs[18][10] ),
    .A3(\regs[19][10] ),
    .S0(_03270_),
    .S1(_03304_),
    .X(_03800_));
 sky130_fd_sc_hd__mux4_1 _09480_ (.A0(\regs[20][10] ),
    .A1(\regs[21][10] ),
    .A2(\regs[22][10] ),
    .A3(\regs[23][10] ),
    .S0(_02280_),
    .S1(_03250_),
    .X(_03801_));
 sky130_fd_sc_hd__or2_1 _09481_ (.A(_03274_),
    .B(_03801_),
    .X(_03802_));
 sky130_fd_sc_hd__o211a_1 _09482_ (.A1(_03357_),
    .A2(_03800_),
    .B1(_03802_),
    .C1(_03258_),
    .X(_03803_));
 sky130_fd_sc_hd__mux4_1 _09483_ (.A0(\regs[12][10] ),
    .A1(\regs[13][10] ),
    .A2(\regs[14][10] ),
    .A3(\regs[15][10] ),
    .S0(_03238_),
    .S1(_03395_),
    .X(_03804_));
 sky130_fd_sc_hd__mux4_1 _09484_ (.A0(\regs[8][10] ),
    .A1(\regs[9][10] ),
    .A2(\regs[10][10] ),
    .A3(\regs[11][10] ),
    .S0(_03400_),
    .S1(_03245_),
    .X(_03805_));
 sky130_fd_sc_hd__or2_1 _09485_ (.A(_02271_),
    .B(_03805_),
    .X(_03806_));
 sky130_fd_sc_hd__o211a_1 _09486_ (.A1(_03236_),
    .A2(_03804_),
    .B1(_03806_),
    .C1(_02267_),
    .X(_03807_));
 sky130_fd_sc_hd__mux4_1 _09487_ (.A0(\regs[0][10] ),
    .A1(\regs[1][10] ),
    .A2(\regs[2][10] ),
    .A3(\regs[3][10] ),
    .S0(_03400_),
    .S1(_03401_),
    .X(_03808_));
 sky130_fd_sc_hd__mux4_1 _09488_ (.A0(\regs[4][10] ),
    .A1(\regs[5][10] ),
    .A2(\regs[6][10] ),
    .A3(\regs[7][10] ),
    .S0(_03237_),
    .S1(_03239_),
    .X(_03809_));
 sky130_fd_sc_hd__mux2_1 _09489_ (.A0(_03808_),
    .A1(_03809_),
    .S(_03254_),
    .X(_03810_));
 sky130_fd_sc_hd__a21o_1 _09490_ (.A1(_03309_),
    .A2(_03810_),
    .B1(net18),
    .X(_03811_));
 sky130_fd_sc_hd__o32a_1 _09491_ (.A1(_02264_),
    .A2(_03799_),
    .A3(_03803_),
    .B1(_03807_),
    .B2(_03811_),
    .X(_03812_));
 sky130_fd_sc_hd__mux2_1 _09492_ (.A0(\rs2_content[10] ),
    .A1(_03812_),
    .S(_02253_),
    .X(_03813_));
 sky130_fd_sc_hd__clkbuf_1 _09493_ (.A(_03813_),
    .X(_01322_));
 sky130_fd_sc_hd__mux4_1 _09494_ (.A0(\regs[12][9] ),
    .A1(\regs[13][9] ),
    .A2(\regs[14][9] ),
    .A3(\regs[15][9] ),
    .S0(_03300_),
    .S1(_03291_),
    .X(_03814_));
 sky130_fd_sc_hd__or2_1 _09495_ (.A(_03362_),
    .B(_03814_),
    .X(_03815_));
 sky130_fd_sc_hd__mux4_1 _09496_ (.A0(\regs[8][9] ),
    .A1(\regs[9][9] ),
    .A2(\regs[10][9] ),
    .A3(\regs[11][9] ),
    .S0(_03554_),
    .S1(_03555_),
    .X(_03816_));
 sky130_fd_sc_hd__o21a_1 _09497_ (.A1(_03316_),
    .A2(_03816_),
    .B1(_03297_),
    .X(_03817_));
 sky130_fd_sc_hd__mux4_1 _09498_ (.A0(\regs[0][9] ),
    .A1(\regs[1][9] ),
    .A2(\regs[2][9] ),
    .A3(\regs[3][9] ),
    .S0(_03303_),
    .S1(_03305_),
    .X(_03818_));
 sky130_fd_sc_hd__mux4_1 _09499_ (.A0(\regs[4][9] ),
    .A1(\regs[5][9] ),
    .A2(\regs[6][9] ),
    .A3(\regs[7][9] ),
    .S0(_03318_),
    .S1(_03336_),
    .X(_03819_));
 sky130_fd_sc_hd__mux2_1 _09500_ (.A0(_03818_),
    .A1(_03819_),
    .S(_03339_),
    .X(_03820_));
 sky130_fd_sc_hd__a22o_1 _09501_ (.A1(_03815_),
    .A2(_03817_),
    .B1(_03820_),
    .B2(_03310_),
    .X(_03821_));
 sky130_fd_sc_hd__mux4_1 _09502_ (.A0(\regs[20][9] ),
    .A1(\regs[21][9] ),
    .A2(\regs[22][9] ),
    .A3(\regs[23][9] ),
    .S0(_03484_),
    .S1(_03485_),
    .X(_03822_));
 sky130_fd_sc_hd__mux4_1 _09503_ (.A0(\regs[16][9] ),
    .A1(\regs[17][9] ),
    .A2(\regs[18][9] ),
    .A3(\regs[19][9] ),
    .S0(_03487_),
    .S1(_03488_),
    .X(_03823_));
 sky130_fd_sc_hd__mux2_1 _09504_ (.A0(_03822_),
    .A1(_03823_),
    .S(_03394_),
    .X(_03824_));
 sky130_fd_sc_hd__mux2_1 _09505_ (.A0(\regs[30][9] ),
    .A1(\regs[31][9] ),
    .S(_03346_),
    .X(_03825_));
 sky130_fd_sc_hd__and2_1 _09506_ (.A(_03341_),
    .B(_03825_),
    .X(_03826_));
 sky130_fd_sc_hd__mux2_1 _09507_ (.A0(\regs[28][9] ),
    .A1(\regs[29][9] ),
    .S(_03327_),
    .X(_03827_));
 sky130_fd_sc_hd__a21o_1 _09508_ (.A1(_03329_),
    .A2(_03827_),
    .B1(_03394_),
    .X(_03828_));
 sky130_fd_sc_hd__or2b_1 _09509_ (.A(\regs[27][9] ),
    .B_N(_03363_),
    .X(_03829_));
 sky130_fd_sc_hd__o21a_1 _09510_ (.A1(_03363_),
    .A2(\regs[26][9] ),
    .B1(_03262_),
    .X(_03830_));
 sky130_fd_sc_hd__mux2_1 _09511_ (.A0(\regs[24][9] ),
    .A1(\regs[25][9] ),
    .S(_03343_),
    .X(_03831_));
 sky130_fd_sc_hd__a221o_1 _09512_ (.A1(_03829_),
    .A2(_03830_),
    .B1(_03831_),
    .B2(_03356_),
    .C1(_02272_),
    .X(_03832_));
 sky130_fd_sc_hd__o211a_1 _09513_ (.A1(_03826_),
    .A2(_03828_),
    .B1(_03832_),
    .C1(_02268_),
    .X(_03833_));
 sky130_fd_sc_hd__a211o_1 _09514_ (.A1(_03334_),
    .A2(_03824_),
    .B1(_03833_),
    .C1(_03500_),
    .X(_03834_));
 sky130_fd_sc_hd__o221a_1 _09515_ (.A1(\rs2_content[9] ),
    .A2(_02993_),
    .B1(_02265_),
    .B2(_03821_),
    .C1(_03834_),
    .X(_01321_));
 sky130_fd_sc_hd__mux2_1 _09516_ (.A0(\regs[30][8] ),
    .A1(\regs[31][8] ),
    .S(_03386_),
    .X(_03835_));
 sky130_fd_sc_hd__and2_1 _09517_ (.A(_03240_),
    .B(_03835_),
    .X(_03836_));
 sky130_fd_sc_hd__mux2_1 _09518_ (.A0(\regs[28][8] ),
    .A1(\regs[29][8] ),
    .S(_03342_),
    .X(_03837_));
 sky130_fd_sc_hd__a21o_1 _09519_ (.A1(_03355_),
    .A2(_03837_),
    .B1(_03235_),
    .X(_03838_));
 sky130_fd_sc_hd__or2b_1 _09520_ (.A(\regs[27][8] ),
    .B_N(_03384_),
    .X(_03839_));
 sky130_fd_sc_hd__o21a_1 _09521_ (.A1(_03384_),
    .A2(\regs[26][8] ),
    .B1(_03250_),
    .X(_03840_));
 sky130_fd_sc_hd__mux2_1 _09522_ (.A0(\regs[24][8] ),
    .A1(\regs[25][8] ),
    .S(_02281_),
    .X(_03841_));
 sky130_fd_sc_hd__a221o_1 _09523_ (.A1(_03839_),
    .A2(_03840_),
    .B1(_03841_),
    .B2(_03272_),
    .C1(net16),
    .X(_03842_));
 sky130_fd_sc_hd__o211a_1 _09524_ (.A1(_03836_),
    .A2(_03838_),
    .B1(_03842_),
    .C1(_03266_),
    .X(_03843_));
 sky130_fd_sc_hd__mux4_1 _09525_ (.A0(\regs[16][8] ),
    .A1(\regs[17][8] ),
    .A2(\regs[18][8] ),
    .A3(\regs[19][8] ),
    .S0(_03270_),
    .S1(_03304_),
    .X(_03844_));
 sky130_fd_sc_hd__mux4_1 _09526_ (.A0(\regs[20][8] ),
    .A1(\regs[21][8] ),
    .A2(\regs[22][8] ),
    .A3(\regs[23][8] ),
    .S0(_02280_),
    .S1(net15),
    .X(_03845_));
 sky130_fd_sc_hd__or2_1 _09527_ (.A(_03274_),
    .B(_03845_),
    .X(_03846_));
 sky130_fd_sc_hd__o211a_1 _09528_ (.A1(_03357_),
    .A2(_03844_),
    .B1(_03846_),
    .C1(_03258_),
    .X(_03847_));
 sky130_fd_sc_hd__mux4_1 _09529_ (.A0(\regs[12][8] ),
    .A1(\regs[13][8] ),
    .A2(\regs[14][8] ),
    .A3(\regs[15][8] ),
    .S0(_03238_),
    .S1(_03395_),
    .X(_03848_));
 sky130_fd_sc_hd__mux4_1 _09530_ (.A0(\regs[8][8] ),
    .A1(\regs[9][8] ),
    .A2(\regs[10][8] ),
    .A3(\regs[11][8] ),
    .S0(_03400_),
    .S1(_03245_),
    .X(_03849_));
 sky130_fd_sc_hd__or2_1 _09531_ (.A(_02271_),
    .B(_03849_),
    .X(_03850_));
 sky130_fd_sc_hd__o211a_1 _09532_ (.A1(_03236_),
    .A2(_03848_),
    .B1(_03850_),
    .C1(_02267_),
    .X(_03851_));
 sky130_fd_sc_hd__mux4_1 _09533_ (.A0(\regs[0][8] ),
    .A1(\regs[1][8] ),
    .A2(\regs[2][8] ),
    .A3(\regs[3][8] ),
    .S0(_03400_),
    .S1(_03401_),
    .X(_03852_));
 sky130_fd_sc_hd__mux4_1 _09534_ (.A0(\regs[4][8] ),
    .A1(\regs[5][8] ),
    .A2(\regs[6][8] ),
    .A3(\regs[7][8] ),
    .S0(_03237_),
    .S1(_03239_),
    .X(_03853_));
 sky130_fd_sc_hd__mux2_1 _09535_ (.A0(_03852_),
    .A1(_03853_),
    .S(_03254_),
    .X(_03854_));
 sky130_fd_sc_hd__a21o_1 _09536_ (.A1(_03309_),
    .A2(_03854_),
    .B1(net18),
    .X(_03855_));
 sky130_fd_sc_hd__o32a_1 _09537_ (.A1(_02263_),
    .A2(_03843_),
    .A3(_03847_),
    .B1(_03851_),
    .B2(_03855_),
    .X(_03856_));
 sky130_fd_sc_hd__mux2_1 _09538_ (.A0(\rs2_content[8] ),
    .A1(_03856_),
    .S(_02253_),
    .X(_03857_));
 sky130_fd_sc_hd__clkbuf_1 _09539_ (.A(_03857_),
    .X(_01320_));
 sky130_fd_sc_hd__mux4_1 _09540_ (.A0(\regs[0][7] ),
    .A1(\regs[1][7] ),
    .A2(\regs[2][7] ),
    .A3(\regs[3][7] ),
    .S0(_03550_),
    .S1(_03551_),
    .X(_03858_));
 sky130_fd_sc_hd__mux4_1 _09541_ (.A0(\regs[4][7] ),
    .A1(\regs[5][7] ),
    .A2(\regs[6][7] ),
    .A3(\regs[7][7] ),
    .S0(_03370_),
    .S1(_03371_),
    .X(_03859_));
 sky130_fd_sc_hd__mux2_1 _09542_ (.A0(_03858_),
    .A1(_03859_),
    .S(_03374_),
    .X(_03860_));
 sky130_fd_sc_hd__mux4_1 _09543_ (.A0(\regs[12][7] ),
    .A1(\regs[13][7] ),
    .A2(\regs[14][7] ),
    .A3(\regs[15][7] ),
    .S0(_03554_),
    .S1(_03555_),
    .X(_03861_));
 sky130_fd_sc_hd__or2_1 _09544_ (.A(_03288_),
    .B(_03861_),
    .X(_03862_));
 sky130_fd_sc_hd__mux4_1 _09545_ (.A0(\regs[8][7] ),
    .A1(\regs[9][7] ),
    .A2(\regs[10][7] ),
    .A3(\regs[11][7] ),
    .S0(_03534_),
    .S1(_03295_),
    .X(_03863_));
 sky130_fd_sc_hd__o21a_1 _09546_ (.A1(_02273_),
    .A2(_03863_),
    .B1(_03359_),
    .X(_03864_));
 sky130_fd_sc_hd__a22o_1 _09547_ (.A1(_03376_),
    .A2(_03860_),
    .B1(_03862_),
    .B2(_03864_),
    .X(_03865_));
 sky130_fd_sc_hd__mux4_1 _09548_ (.A0(\regs[16][7] ),
    .A1(\regs[17][7] ),
    .A2(\regs[18][7] ),
    .A3(\regs[19][7] ),
    .S0(_03484_),
    .S1(_03485_),
    .X(_03866_));
 sky130_fd_sc_hd__mux4_1 _09549_ (.A0(\regs[20][7] ),
    .A1(\regs[21][7] ),
    .A2(\regs[22][7] ),
    .A3(\regs[23][7] ),
    .S0(_03487_),
    .S1(_03488_),
    .X(_03867_));
 sky130_fd_sc_hd__mux2_1 _09550_ (.A0(_03866_),
    .A1(_03867_),
    .S(_03307_),
    .X(_03868_));
 sky130_fd_sc_hd__mux2_1 _09551_ (.A0(\regs[30][7] ),
    .A1(\regs[31][7] ),
    .S(_03327_),
    .X(_03869_));
 sky130_fd_sc_hd__mux2_1 _09552_ (.A0(\regs[28][7] ),
    .A1(\regs[29][7] ),
    .S(_03349_),
    .X(_03870_));
 sky130_fd_sc_hd__a21o_1 _09553_ (.A1(_03543_),
    .A2(_03870_),
    .B1(_03566_),
    .X(_03871_));
 sky130_fd_sc_hd__a21o_1 _09554_ (.A1(_03341_),
    .A2(_03869_),
    .B1(_03871_),
    .X(_03872_));
 sky130_fd_sc_hd__or2b_1 _09555_ (.A(\regs[27][7] ),
    .B_N(_03569_),
    .X(_03873_));
 sky130_fd_sc_hd__o21a_1 _09556_ (.A1(_03539_),
    .A2(\regs[26][7] ),
    .B1(_03352_),
    .X(_03874_));
 sky130_fd_sc_hd__mux2_1 _09557_ (.A0(\regs[24][7] ),
    .A1(\regs[25][7] ),
    .S(_03261_),
    .X(_03875_));
 sky130_fd_sc_hd__a221o_1 _09558_ (.A1(_03873_),
    .A2(_03874_),
    .B1(_03875_),
    .B2(_03320_),
    .C1(_03255_),
    .X(_03876_));
 sky130_fd_sc_hd__and3_1 _09559_ (.A(_03368_),
    .B(_03872_),
    .C(_03876_),
    .X(_03877_));
 sky130_fd_sc_hd__a211o_1 _09560_ (.A1(_03334_),
    .A2(_03868_),
    .B1(_03877_),
    .C1(_03500_),
    .X(_03878_));
 sky130_fd_sc_hd__o221a_1 _09561_ (.A1(\rs2_content[7] ),
    .A2(_02993_),
    .B1(_02265_),
    .B2(_03865_),
    .C1(_03878_),
    .X(_01319_));
 sky130_fd_sc_hd__mux4_1 _09562_ (.A0(\regs[0][6] ),
    .A1(\regs[1][6] ),
    .A2(\regs[2][6] ),
    .A3(\regs[3][6] ),
    .S0(_03550_),
    .S1(_03551_),
    .X(_03879_));
 sky130_fd_sc_hd__mux4_1 _09563_ (.A0(\regs[4][6] ),
    .A1(\regs[5][6] ),
    .A2(\regs[6][6] ),
    .A3(\regs[7][6] ),
    .S0(_03370_),
    .S1(_03371_),
    .X(_03880_));
 sky130_fd_sc_hd__mux2_1 _09564_ (.A0(_03879_),
    .A1(_03880_),
    .S(_03374_),
    .X(_03881_));
 sky130_fd_sc_hd__mux4_1 _09565_ (.A0(\regs[12][6] ),
    .A1(\regs[13][6] ),
    .A2(\regs[14][6] ),
    .A3(\regs[15][6] ),
    .S0(_03554_),
    .S1(_03555_),
    .X(_03882_));
 sky130_fd_sc_hd__or2_1 _09566_ (.A(_03288_),
    .B(_03882_),
    .X(_03883_));
 sky130_fd_sc_hd__mux4_1 _09567_ (.A0(\regs[8][6] ),
    .A1(\regs[9][6] ),
    .A2(\regs[10][6] ),
    .A3(\regs[11][6] ),
    .S0(_03294_),
    .S1(_03295_),
    .X(_03884_));
 sky130_fd_sc_hd__o21a_1 _09568_ (.A1(_02273_),
    .A2(_03884_),
    .B1(_03359_),
    .X(_03885_));
 sky130_fd_sc_hd__a22o_1 _09569_ (.A1(_03376_),
    .A2(_03881_),
    .B1(_03883_),
    .B2(_03885_),
    .X(_03886_));
 sky130_fd_sc_hd__mux4_1 _09570_ (.A0(\regs[16][6] ),
    .A1(\regs[17][6] ),
    .A2(\regs[18][6] ),
    .A3(\regs[19][6] ),
    .S0(_03484_),
    .S1(_03485_),
    .X(_03887_));
 sky130_fd_sc_hd__mux4_1 _09571_ (.A0(\regs[20][6] ),
    .A1(\regs[21][6] ),
    .A2(\regs[22][6] ),
    .A3(\regs[23][6] ),
    .S0(_03487_),
    .S1(_03488_),
    .X(_03888_));
 sky130_fd_sc_hd__mux2_1 _09572_ (.A0(_03887_),
    .A1(_03888_),
    .S(_03307_),
    .X(_03889_));
 sky130_fd_sc_hd__mux2_1 _09573_ (.A0(\regs[30][6] ),
    .A1(\regs[31][6] ),
    .S(_03346_),
    .X(_03890_));
 sky130_fd_sc_hd__mux2_1 _09574_ (.A0(\regs[28][6] ),
    .A1(\regs[29][6] ),
    .S(_03349_),
    .X(_03891_));
 sky130_fd_sc_hd__a21o_1 _09575_ (.A1(_03543_),
    .A2(_03891_),
    .B1(_03566_),
    .X(_03892_));
 sky130_fd_sc_hd__a21o_1 _09576_ (.A1(_03341_),
    .A2(_03890_),
    .B1(_03892_),
    .X(_03893_));
 sky130_fd_sc_hd__or2b_1 _09577_ (.A(\regs[27][6] ),
    .B_N(_03569_),
    .X(_03894_));
 sky130_fd_sc_hd__o21a_1 _09578_ (.A1(_03539_),
    .A2(\regs[26][6] ),
    .B1(_03395_),
    .X(_03895_));
 sky130_fd_sc_hd__mux2_1 _09579_ (.A0(\regs[24][6] ),
    .A1(\regs[25][6] ),
    .S(_03261_),
    .X(_03896_));
 sky130_fd_sc_hd__a221o_1 _09580_ (.A1(_03894_),
    .A2(_03895_),
    .B1(_03896_),
    .B2(_03320_),
    .C1(_03255_),
    .X(_03897_));
 sky130_fd_sc_hd__and3_1 _09581_ (.A(_03368_),
    .B(_03893_),
    .C(_03897_),
    .X(_03898_));
 sky130_fd_sc_hd__a211o_1 _09582_ (.A1(_03334_),
    .A2(_03889_),
    .B1(_03898_),
    .C1(_03500_),
    .X(_03899_));
 sky130_fd_sc_hd__o221a_1 _09583_ (.A1(\rs2_content[6] ),
    .A2(_02993_),
    .B1(_02265_),
    .B2(_03886_),
    .C1(_03899_),
    .X(_01318_));
 sky130_fd_sc_hd__mux4_1 _09584_ (.A0(\regs[12][5] ),
    .A1(\regs[13][5] ),
    .A2(\regs[14][5] ),
    .A3(\regs[15][5] ),
    .S0(_03249_),
    .S1(_03240_),
    .X(_03900_));
 sky130_fd_sc_hd__or2_1 _09585_ (.A(_03287_),
    .B(_03900_),
    .X(_03901_));
 sky130_fd_sc_hd__mux4_1 _09586_ (.A0(\regs[8][5] ),
    .A1(\regs[9][5] ),
    .A2(\regs[10][5] ),
    .A3(\regs[11][5] ),
    .S0(_03238_),
    .S1(_03246_),
    .X(_03902_));
 sky130_fd_sc_hd__o21a_1 _09587_ (.A1(_03244_),
    .A2(_03902_),
    .B1(_02267_),
    .X(_03903_));
 sky130_fd_sc_hd__mux4_1 _09588_ (.A0(\regs[0][5] ),
    .A1(\regs[1][5] ),
    .A2(\regs[2][5] ),
    .A3(\regs[3][5] ),
    .S0(_03249_),
    .S1(_03251_),
    .X(_03904_));
 sky130_fd_sc_hd__mux4_1 _09589_ (.A0(\regs[4][5] ),
    .A1(\regs[5][5] ),
    .A2(\regs[6][5] ),
    .A3(\regs[7][5] ),
    .S0(_03277_),
    .S1(_03251_),
    .X(_03905_));
 sky130_fd_sc_hd__mux2_1 _09590_ (.A0(_03904_),
    .A1(_03905_),
    .S(_03243_),
    .X(_03906_));
 sky130_fd_sc_hd__a22o_1 _09591_ (.A1(_03901_),
    .A2(_03903_),
    .B1(_03906_),
    .B2(_03309_),
    .X(_03907_));
 sky130_fd_sc_hd__mux4_1 _09592_ (.A0(\regs[16][5] ),
    .A1(\regs[17][5] ),
    .A2(\regs[18][5] ),
    .A3(\regs[19][5] ),
    .S0(_02282_),
    .S1(_03262_),
    .X(_03908_));
 sky130_fd_sc_hd__mux4_1 _09593_ (.A0(\regs[20][5] ),
    .A1(\regs[21][5] ),
    .A2(\regs[22][5] ),
    .A3(\regs[23][5] ),
    .S0(_02282_),
    .S1(_03352_),
    .X(_03909_));
 sky130_fd_sc_hd__mux2_1 _09594_ (.A0(_03908_),
    .A1(_03909_),
    .S(_02272_),
    .X(_03910_));
 sky130_fd_sc_hd__mux2_1 _09595_ (.A0(\regs[30][5] ),
    .A1(\regs[31][5] ),
    .S(_03299_),
    .X(_03911_));
 sky130_fd_sc_hd__mux2_1 _09596_ (.A0(\regs[28][5] ),
    .A1(\regs[29][5] ),
    .S(_03269_),
    .X(_03912_));
 sky130_fd_sc_hd__a21o_1 _09597_ (.A1(_03272_),
    .A2(_03912_),
    .B1(_03274_),
    .X(_03913_));
 sky130_fd_sc_hd__a21o_1 _09598_ (.A1(_03268_),
    .A2(_03911_),
    .B1(_03913_),
    .X(_03914_));
 sky130_fd_sc_hd__or2b_1 _09599_ (.A(\regs[27][5] ),
    .B_N(_03277_),
    .X(_03915_));
 sky130_fd_sc_hd__o21a_1 _09600_ (.A1(_03289_),
    .A2(\regs[26][5] ),
    .B1(_02276_),
    .X(_03916_));
 sky130_fd_sc_hd__mux2_1 _09601_ (.A0(\regs[24][5] ),
    .A1(\regs[25][5] ),
    .S(_03280_),
    .X(_03917_));
 sky130_fd_sc_hd__a221o_1 _09602_ (.A1(_03915_),
    .A2(_03916_),
    .B1(_03917_),
    .B2(_03282_),
    .C1(_03243_),
    .X(_03918_));
 sky130_fd_sc_hd__a31o_1 _09603_ (.A1(_03267_),
    .A2(_03914_),
    .A3(_03918_),
    .B1(_02263_),
    .X(_03919_));
 sky130_fd_sc_hd__a21o_1 _09604_ (.A1(_03259_),
    .A2(_03910_),
    .B1(_03919_),
    .X(_03920_));
 sky130_fd_sc_hd__o211a_1 _09605_ (.A1(_03233_),
    .A2(_03907_),
    .B1(_03920_),
    .C1(_02254_),
    .X(_03921_));
 sky130_fd_sc_hd__a21o_1 _09606_ (.A1(\rs2_content[5] ),
    .A2(_02543_),
    .B1(_03921_),
    .X(_01317_));
 sky130_fd_sc_hd__mux4_1 _09607_ (.A0(\regs[4][4] ),
    .A1(\regs[5][4] ),
    .A2(\regs[6][4] ),
    .A3(\regs[7][4] ),
    .S0(_03550_),
    .S1(_03551_),
    .X(_03922_));
 sky130_fd_sc_hd__mux4_1 _09608_ (.A0(\regs[0][4] ),
    .A1(\regs[1][4] ),
    .A2(\regs[2][4] ),
    .A3(\regs[3][4] ),
    .S0(_03370_),
    .S1(_03371_),
    .X(_03923_));
 sky130_fd_sc_hd__mux2_1 _09609_ (.A0(_03922_),
    .A1(_03923_),
    .S(_03394_),
    .X(_03924_));
 sky130_fd_sc_hd__mux4_1 _09610_ (.A0(\regs[12][4] ),
    .A1(\regs[13][4] ),
    .A2(\regs[14][4] ),
    .A3(\regs[15][4] ),
    .S0(_03554_),
    .S1(_03555_),
    .X(_03925_));
 sky130_fd_sc_hd__or2_1 _09611_ (.A(_03288_),
    .B(_03925_),
    .X(_03926_));
 sky130_fd_sc_hd__mux4_1 _09612_ (.A0(\regs[8][4] ),
    .A1(\regs[9][4] ),
    .A2(\regs[10][4] ),
    .A3(\regs[11][4] ),
    .S0(_03294_),
    .S1(_03295_),
    .X(_03927_));
 sky130_fd_sc_hd__o21a_1 _09613_ (.A1(_02273_),
    .A2(_03927_),
    .B1(_03359_),
    .X(_03928_));
 sky130_fd_sc_hd__a22o_1 _09614_ (.A1(_03376_),
    .A2(_03924_),
    .B1(_03926_),
    .B2(_03928_),
    .X(_03929_));
 sky130_fd_sc_hd__mux4_1 _09615_ (.A0(\regs[16][4] ),
    .A1(\regs[17][4] ),
    .A2(\regs[18][4] ),
    .A3(\regs[19][4] ),
    .S0(_03484_),
    .S1(_03485_),
    .X(_03930_));
 sky130_fd_sc_hd__mux4_1 _09616_ (.A0(\regs[20][4] ),
    .A1(\regs[21][4] ),
    .A2(\regs[22][4] ),
    .A3(\regs[23][4] ),
    .S0(_03487_),
    .S1(_03488_),
    .X(_03931_));
 sky130_fd_sc_hd__mux2_1 _09617_ (.A0(_03930_),
    .A1(_03931_),
    .S(_03307_),
    .X(_03932_));
 sky130_fd_sc_hd__mux2_1 _09618_ (.A0(\regs[30][4] ),
    .A1(\regs[31][4] ),
    .S(_03346_),
    .X(_03933_));
 sky130_fd_sc_hd__mux2_1 _09619_ (.A0(\regs[28][4] ),
    .A1(\regs[29][4] ),
    .S(_03349_),
    .X(_03934_));
 sky130_fd_sc_hd__a21o_1 _09620_ (.A1(_03282_),
    .A2(_03934_),
    .B1(_03566_),
    .X(_03935_));
 sky130_fd_sc_hd__a21o_1 _09621_ (.A1(_03341_),
    .A2(_03933_),
    .B1(_03935_),
    .X(_03936_));
 sky130_fd_sc_hd__or2b_1 _09622_ (.A(\regs[27][4] ),
    .B_N(_03569_),
    .X(_03937_));
 sky130_fd_sc_hd__o21a_1 _09623_ (.A1(_03539_),
    .A2(\regs[26][4] ),
    .B1(_03395_),
    .X(_03938_));
 sky130_fd_sc_hd__mux2_1 _09624_ (.A0(\regs[24][4] ),
    .A1(\regs[25][4] ),
    .S(_03261_),
    .X(_03939_));
 sky130_fd_sc_hd__a221o_1 _09625_ (.A1(_03937_),
    .A2(_03938_),
    .B1(_03939_),
    .B2(_03320_),
    .C1(_03255_),
    .X(_03940_));
 sky130_fd_sc_hd__and3_1 _09626_ (.A(_03368_),
    .B(_03936_),
    .C(_03940_),
    .X(_03941_));
 sky130_fd_sc_hd__a211o_1 _09627_ (.A1(_03334_),
    .A2(_03932_),
    .B1(_03941_),
    .C1(_03500_),
    .X(_03942_));
 sky130_fd_sc_hd__o221a_1 _09628_ (.A1(\rs2_content[4] ),
    .A2(_02993_),
    .B1(_02265_),
    .B2(_03929_),
    .C1(_03942_),
    .X(_01316_));
 sky130_fd_sc_hd__mux2_1 _09629_ (.A0(\regs[30][3] ),
    .A1(\regs[31][3] ),
    .S(_03386_),
    .X(_03943_));
 sky130_fd_sc_hd__and2_1 _09630_ (.A(_03240_),
    .B(_03943_),
    .X(_03944_));
 sky130_fd_sc_hd__mux2_1 _09631_ (.A0(\regs[28][3] ),
    .A1(\regs[29][3] ),
    .S(_03342_),
    .X(_03945_));
 sky130_fd_sc_hd__a21o_1 _09632_ (.A1(_03355_),
    .A2(_03945_),
    .B1(_03235_),
    .X(_03946_));
 sky130_fd_sc_hd__or2b_1 _09633_ (.A(\regs[27][3] ),
    .B_N(_03384_),
    .X(_03947_));
 sky130_fd_sc_hd__o21a_1 _09634_ (.A1(_03384_),
    .A2(\regs[26][3] ),
    .B1(_03250_),
    .X(_03948_));
 sky130_fd_sc_hd__mux2_1 _09635_ (.A0(\regs[24][3] ),
    .A1(\regs[25][3] ),
    .S(_02281_),
    .X(_03949_));
 sky130_fd_sc_hd__a221o_1 _09636_ (.A1(_03947_),
    .A2(_03948_),
    .B1(_03949_),
    .B2(_03272_),
    .C1(net16),
    .X(_03950_));
 sky130_fd_sc_hd__o211a_1 _09637_ (.A1(_03944_),
    .A2(_03946_),
    .B1(_03950_),
    .C1(_03266_),
    .X(_03951_));
 sky130_fd_sc_hd__mux4_1 _09638_ (.A0(\regs[16][3] ),
    .A1(\regs[17][3] ),
    .A2(\regs[18][3] ),
    .A3(\regs[19][3] ),
    .S0(_03270_),
    .S1(_03304_),
    .X(_03952_));
 sky130_fd_sc_hd__mux4_1 _09639_ (.A0(\regs[20][3] ),
    .A1(\regs[21][3] ),
    .A2(\regs[22][3] ),
    .A3(\regs[23][3] ),
    .S0(_02280_),
    .S1(net15),
    .X(_03953_));
 sky130_fd_sc_hd__or2_1 _09640_ (.A(_03274_),
    .B(_03953_),
    .X(_03954_));
 sky130_fd_sc_hd__o211a_1 _09641_ (.A1(_03357_),
    .A2(_03952_),
    .B1(_03954_),
    .C1(_03258_),
    .X(_03955_));
 sky130_fd_sc_hd__mux4_1 _09642_ (.A0(\regs[12][3] ),
    .A1(\regs[13][3] ),
    .A2(\regs[14][3] ),
    .A3(\regs[15][3] ),
    .S0(_03238_),
    .S1(_03395_),
    .X(_03956_));
 sky130_fd_sc_hd__mux4_1 _09643_ (.A0(\regs[8][3] ),
    .A1(\regs[9][3] ),
    .A2(\regs[10][3] ),
    .A3(\regs[11][3] ),
    .S0(_03400_),
    .S1(_03245_),
    .X(_03957_));
 sky130_fd_sc_hd__or2_1 _09644_ (.A(_02271_),
    .B(_03957_),
    .X(_03958_));
 sky130_fd_sc_hd__o211a_1 _09645_ (.A1(_03236_),
    .A2(_03956_),
    .B1(_03958_),
    .C1(_02267_),
    .X(_03959_));
 sky130_fd_sc_hd__mux4_1 _09646_ (.A0(\regs[0][3] ),
    .A1(\regs[1][3] ),
    .A2(\regs[2][3] ),
    .A3(\regs[3][3] ),
    .S0(_03400_),
    .S1(_03401_),
    .X(_03960_));
 sky130_fd_sc_hd__mux4_1 _09647_ (.A0(\regs[4][3] ),
    .A1(\regs[5][3] ),
    .A2(\regs[6][3] ),
    .A3(\regs[7][3] ),
    .S0(_03237_),
    .S1(_03239_),
    .X(_03961_));
 sky130_fd_sc_hd__mux2_1 _09648_ (.A0(_03960_),
    .A1(_03961_),
    .S(_03254_),
    .X(_03962_));
 sky130_fd_sc_hd__a21o_1 _09649_ (.A1(_03258_),
    .A2(_03962_),
    .B1(net18),
    .X(_03963_));
 sky130_fd_sc_hd__o32a_2 _09650_ (.A1(_02263_),
    .A2(_03951_),
    .A3(_03955_),
    .B1(_03959_),
    .B2(_03963_),
    .X(_03964_));
 sky130_fd_sc_hd__mux2_1 _09651_ (.A0(_01770_),
    .A1(_03964_),
    .S(_02253_),
    .X(_03965_));
 sky130_fd_sc_hd__clkbuf_1 _09652_ (.A(_03965_),
    .X(_01315_));
 sky130_fd_sc_hd__mux4_1 _09653_ (.A0(\regs[0][2] ),
    .A1(\regs[1][2] ),
    .A2(\regs[2][2] ),
    .A3(\regs[3][2] ),
    .S0(_03550_),
    .S1(_03551_),
    .X(_03966_));
 sky130_fd_sc_hd__mux4_1 _09654_ (.A0(\regs[4][2] ),
    .A1(\regs[5][2] ),
    .A2(\regs[6][2] ),
    .A3(\regs[7][2] ),
    .S0(_03370_),
    .S1(_03371_),
    .X(_03967_));
 sky130_fd_sc_hd__mux2_1 _09655_ (.A0(_03966_),
    .A1(_03967_),
    .S(_03374_),
    .X(_03968_));
 sky130_fd_sc_hd__mux4_1 _09656_ (.A0(\regs[12][2] ),
    .A1(\regs[13][2] ),
    .A2(\regs[14][2] ),
    .A3(\regs[15][2] ),
    .S0(_03554_),
    .S1(_03485_),
    .X(_03969_));
 sky130_fd_sc_hd__or2_1 _09657_ (.A(_03288_),
    .B(_03969_),
    .X(_03970_));
 sky130_fd_sc_hd__mux4_1 _09658_ (.A0(\regs[8][2] ),
    .A1(\regs[9][2] ),
    .A2(\regs[10][2] ),
    .A3(\regs[11][2] ),
    .S0(_03294_),
    .S1(_03295_),
    .X(_03971_));
 sky130_fd_sc_hd__o21a_1 _09659_ (.A1(_02273_),
    .A2(_03971_),
    .B1(_03359_),
    .X(_03972_));
 sky130_fd_sc_hd__a22o_1 _09660_ (.A1(_03376_),
    .A2(_03968_),
    .B1(_03970_),
    .B2(_03972_),
    .X(_03973_));
 sky130_fd_sc_hd__mux4_1 _09661_ (.A0(\regs[16][2] ),
    .A1(\regs[17][2] ),
    .A2(\regs[18][2] ),
    .A3(\regs[19][2] ),
    .S0(_03484_),
    .S1(_03488_),
    .X(_03974_));
 sky130_fd_sc_hd__mux4_1 _09662_ (.A0(\regs[20][2] ),
    .A1(\regs[21][2] ),
    .A2(\regs[22][2] ),
    .A3(\regs[23][2] ),
    .S0(_03487_),
    .S1(_03291_),
    .X(_03975_));
 sky130_fd_sc_hd__mux2_1 _09663_ (.A0(_03974_),
    .A1(_03975_),
    .S(_03307_),
    .X(_03976_));
 sky130_fd_sc_hd__mux2_1 _09664_ (.A0(\regs[30][2] ),
    .A1(\regs[31][2] ),
    .S(_03346_),
    .X(_03977_));
 sky130_fd_sc_hd__mux2_1 _09665_ (.A0(\regs[28][2] ),
    .A1(\regs[29][2] ),
    .S(_03280_),
    .X(_03978_));
 sky130_fd_sc_hd__a21o_1 _09666_ (.A1(_03282_),
    .A2(_03978_),
    .B1(_03566_),
    .X(_03979_));
 sky130_fd_sc_hd__a21o_1 _09667_ (.A1(_03341_),
    .A2(_03977_),
    .B1(_03979_),
    .X(_03980_));
 sky130_fd_sc_hd__or2b_1 _09668_ (.A(\regs[27][2] ),
    .B_N(_03569_),
    .X(_03981_));
 sky130_fd_sc_hd__o21a_1 _09669_ (.A1(_03539_),
    .A2(\regs[26][2] ),
    .B1(_03395_),
    .X(_03982_));
 sky130_fd_sc_hd__mux2_1 _09670_ (.A0(\regs[24][2] ),
    .A1(\regs[25][2] ),
    .S(_03261_),
    .X(_03983_));
 sky130_fd_sc_hd__a221o_1 _09671_ (.A1(_03981_),
    .A2(_03982_),
    .B1(_03983_),
    .B2(_03320_),
    .C1(_03255_),
    .X(_03984_));
 sky130_fd_sc_hd__and3_1 _09672_ (.A(_03368_),
    .B(_03980_),
    .C(_03984_),
    .X(_03985_));
 sky130_fd_sc_hd__a211o_1 _09673_ (.A1(_03334_),
    .A2(_03976_),
    .B1(_03985_),
    .C1(_03500_),
    .X(_03986_));
 sky130_fd_sc_hd__o221a_2 _09674_ (.A1(_01772_),
    .A2(_02993_),
    .B1(_02265_),
    .B2(_03973_),
    .C1(_03986_),
    .X(_01314_));
 sky130_fd_sc_hd__mux4_1 _09675_ (.A0(\regs[16][1] ),
    .A1(\regs[17][1] ),
    .A2(\regs[18][1] ),
    .A3(\regs[19][1] ),
    .S0(_03335_),
    .S1(_03336_),
    .X(_03987_));
 sky130_fd_sc_hd__mux4_1 _09676_ (.A0(\regs[20][1] ),
    .A1(\regs[21][1] ),
    .A2(\regs[22][1] ),
    .A3(\regs[23][1] ),
    .S0(_03335_),
    .S1(_03336_),
    .X(_03988_));
 sky130_fd_sc_hd__mux2_1 _09677_ (.A0(_03987_),
    .A1(_03988_),
    .S(_03339_),
    .X(_03989_));
 sky130_fd_sc_hd__mux2_1 _09678_ (.A0(\regs[30][1] ),
    .A1(\regs[31][1] ),
    .S(_03343_),
    .X(_03990_));
 sky130_fd_sc_hd__and2_1 _09679_ (.A(_03313_),
    .B(_03990_),
    .X(_03991_));
 sky130_fd_sc_hd__mux2_1 _09680_ (.A0(\regs[28][1] ),
    .A1(\regs[29][1] ),
    .S(_03346_),
    .X(_03992_));
 sky130_fd_sc_hd__a21o_1 _09681_ (.A1(_03356_),
    .A2(_03992_),
    .B1(_03236_),
    .X(_03993_));
 sky130_fd_sc_hd__or2b_1 _09682_ (.A(\regs[27][1] ),
    .B_N(_03350_),
    .X(_03994_));
 sky130_fd_sc_hd__o21a_1 _09683_ (.A1(_03350_),
    .A2(\regs[26][1] ),
    .B1(_03352_),
    .X(_03995_));
 sky130_fd_sc_hd__mux2_1 _09684_ (.A0(\regs[24][1] ),
    .A1(\regs[25][1] ),
    .S(_03343_),
    .X(_03996_));
 sky130_fd_sc_hd__a221o_1 _09685_ (.A1(_03994_),
    .A2(_03995_),
    .B1(_03996_),
    .B2(_03356_),
    .C1(_03357_),
    .X(_03997_));
 sky130_fd_sc_hd__o211a_1 _09686_ (.A1(_03991_),
    .A2(_03993_),
    .B1(_03997_),
    .C1(_03297_),
    .X(_03998_));
 sky130_fd_sc_hd__a211o_1 _09687_ (.A1(_03310_),
    .A2(_03989_),
    .B1(_03998_),
    .C1(_02264_),
    .X(_03999_));
 sky130_fd_sc_hd__mux4_1 _09688_ (.A0(\regs[12][1] ),
    .A1(\regs[13][1] ),
    .A2(\regs[14][1] ),
    .A3(\regs[15][1] ),
    .S0(_03363_),
    .S1(_03268_),
    .X(_04000_));
 sky130_fd_sc_hd__or2_1 _09689_ (.A(_03394_),
    .B(_04000_),
    .X(_04001_));
 sky130_fd_sc_hd__mux4_1 _09690_ (.A0(\regs[8][1] ),
    .A1(\regs[9][1] ),
    .A2(\regs[10][1] ),
    .A3(\regs[11][1] ),
    .S0(_03300_),
    .S1(_03301_),
    .X(_04002_));
 sky130_fd_sc_hd__o21a_1 _09691_ (.A1(_03366_),
    .A2(_04002_),
    .B1(_03267_),
    .X(_04003_));
 sky130_fd_sc_hd__mux4_1 _09692_ (.A0(\regs[0][1] ),
    .A1(\regs[1][1] ),
    .A2(\regs[2][1] ),
    .A3(\regs[3][1] ),
    .S0(_03370_),
    .S1(_03371_),
    .X(_04004_));
 sky130_fd_sc_hd__mux4_1 _09693_ (.A0(\regs[4][1] ),
    .A1(\regs[5][1] ),
    .A2(\regs[6][1] ),
    .A3(\regs[7][1] ),
    .S0(_03350_),
    .S1(_02277_),
    .X(_04005_));
 sky130_fd_sc_hd__mux2_1 _09694_ (.A0(_04004_),
    .A1(_04005_),
    .S(_03374_),
    .X(_04006_));
 sky130_fd_sc_hd__a221o_1 _09695_ (.A1(_04001_),
    .A2(_04003_),
    .B1(_04006_),
    .B2(_03259_),
    .C1(_03233_),
    .X(_04007_));
 sky130_fd_sc_hd__nor2_1 _09696_ (.A(_01779_),
    .B(_02254_),
    .Y(_04008_));
 sky130_fd_sc_hd__a31o_1 _09697_ (.A1(_00001_),
    .A2(_03999_),
    .A3(_04007_),
    .B1(_04008_),
    .X(_01313_));
 sky130_fd_sc_hd__mux4_1 _09698_ (.A0(\regs[12][0] ),
    .A1(\regs[13][0] ),
    .A2(\regs[14][0] ),
    .A3(\regs[15][0] ),
    .S0(_03300_),
    .S1(_03291_),
    .X(_04009_));
 sky130_fd_sc_hd__or2_1 _09699_ (.A(_03362_),
    .B(_04009_),
    .X(_04010_));
 sky130_fd_sc_hd__mux4_1 _09700_ (.A0(\regs[8][0] ),
    .A1(\regs[9][0] ),
    .A2(\regs[10][0] ),
    .A3(\regs[11][0] ),
    .S0(_03554_),
    .S1(_03555_),
    .X(_04011_));
 sky130_fd_sc_hd__o21a_1 _09701_ (.A1(_03316_),
    .A2(_04011_),
    .B1(_03368_),
    .X(_04012_));
 sky130_fd_sc_hd__mux4_1 _09702_ (.A0(\regs[0][0] ),
    .A1(\regs[1][0] ),
    .A2(\regs[2][0] ),
    .A3(\regs[3][0] ),
    .S0(_03303_),
    .S1(_03305_),
    .X(_04013_));
 sky130_fd_sc_hd__mux4_1 _09703_ (.A0(\regs[4][0] ),
    .A1(\regs[5][0] ),
    .A2(\regs[6][0] ),
    .A3(\regs[7][0] ),
    .S0(_03318_),
    .S1(_03336_),
    .X(_04014_));
 sky130_fd_sc_hd__mux2_1 _09704_ (.A0(_04013_),
    .A1(_04014_),
    .S(_03339_),
    .X(_04015_));
 sky130_fd_sc_hd__a22o_1 _09705_ (.A1(_04010_),
    .A2(_04012_),
    .B1(_04015_),
    .B2(_03310_),
    .X(_04016_));
 sky130_fd_sc_hd__mux4_1 _09706_ (.A0(\regs[20][0] ),
    .A1(\regs[21][0] ),
    .A2(\regs[22][0] ),
    .A3(\regs[23][0] ),
    .S0(_02283_),
    .S1(_03313_),
    .X(_04017_));
 sky130_fd_sc_hd__mux4_1 _09707_ (.A0(\regs[16][0] ),
    .A1(\regs[17][0] ),
    .A2(\regs[18][0] ),
    .A3(\regs[19][0] ),
    .S0(_03534_),
    .S1(_03418_),
    .X(_04018_));
 sky130_fd_sc_hd__mux2_1 _09708_ (.A0(_04017_),
    .A1(_04018_),
    .S(_03288_),
    .X(_04019_));
 sky130_fd_sc_hd__or2b_1 _09709_ (.A(\regs[27][0] ),
    .B_N(_03324_),
    .X(_04020_));
 sky130_fd_sc_hd__o21a_1 _09710_ (.A1(_03324_),
    .A2(\regs[26][0] ),
    .B1(_02277_),
    .X(_04021_));
 sky130_fd_sc_hd__mux2_1 _09711_ (.A0(\regs[24][0] ),
    .A1(\regs[25][0] ),
    .S(_03539_),
    .X(_04022_));
 sky130_fd_sc_hd__a221o_1 _09712_ (.A1(_04020_),
    .A2(_04021_),
    .B1(_04022_),
    .B2(_03329_),
    .C1(_03244_),
    .X(_04023_));
 sky130_fd_sc_hd__mux2_1 _09713_ (.A0(\regs[30][0] ),
    .A1(\regs[31][0] ),
    .S(_03335_),
    .X(_04024_));
 sky130_fd_sc_hd__mux2_1 _09714_ (.A0(\regs[28][0] ),
    .A1(\regs[29][0] ),
    .S(_03270_),
    .X(_04025_));
 sky130_fd_sc_hd__a21o_1 _09715_ (.A1(_03543_),
    .A2(_04025_),
    .B1(_03566_),
    .X(_04026_));
 sky130_fd_sc_hd__a21o_1 _09716_ (.A1(_02278_),
    .A2(_04024_),
    .B1(_04026_),
    .X(_04027_));
 sky130_fd_sc_hd__a31o_1 _09717_ (.A1(_02268_),
    .A2(_04023_),
    .A3(_04027_),
    .B1(_03331_),
    .X(_04028_));
 sky130_fd_sc_hd__a21o_1 _09718_ (.A1(_03312_),
    .A2(_04019_),
    .B1(_04028_),
    .X(_04029_));
 sky130_fd_sc_hd__o221a_1 _09719_ (.A1(\rs2_content[0] ),
    .A2(_02993_),
    .B1(_02265_),
    .B2(_04016_),
    .C1(_04029_),
    .X(_01312_));
 sky130_fd_sc_hd__or2_1 _09720_ (.A(_01648_),
    .B(\PC[1] ),
    .X(_04030_));
 sky130_fd_sc_hd__nand2_1 _09721_ (.A(_02275_),
    .B(\PC[1] ),
    .Y(_04031_));
 sky130_fd_sc_hd__or2_1 _09722_ (.A(_02275_),
    .B(\PC[1] ),
    .X(_04032_));
 sky130_fd_sc_hd__xor2_4 _09723_ (.A(_01903_),
    .B(_01904_),
    .X(_04033_));
 sky130_fd_sc_hd__clkbuf_4 _09724_ (.A(_04033_),
    .X(_04034_));
 sky130_fd_sc_hd__a32o_1 _09725_ (.A1(_04031_),
    .A2(_01534_),
    .A3(_04032_),
    .B1(_04034_),
    .B2(_01861_),
    .X(_04035_));
 sky130_fd_sc_hd__a31o_1 _09726_ (.A1(_01649_),
    .A2(_02021_),
    .A3(_04030_),
    .B1(_04035_),
    .X(_04036_));
 sky130_fd_sc_hd__nand2_1 _09727_ (.A(_01985_),
    .B(_01994_),
    .Y(_04037_));
 sky130_fd_sc_hd__mux2_1 _09728_ (.A0(_04036_),
    .A1(\PC[1] ),
    .S(_04037_),
    .X(_04038_));
 sky130_fd_sc_hd__clkbuf_1 _09729_ (.A(_04038_),
    .X(_00831_));
 sky130_fd_sc_hd__o21ai_1 _09730_ (.A1(net1),
    .A2(net34),
    .B1(\core_state[3] ),
    .Y(_04039_));
 sky130_fd_sc_hd__nand2_1 _09731_ (.A(_01529_),
    .B(_04039_),
    .Y(_00003_));
 sky130_fd_sc_hd__a21o_1 _09732_ (.A1(net1),
    .A2(\core_state[2] ),
    .B1(\core_state[0] ),
    .X(_00002_));
 sky130_fd_sc_hd__nor2_1 _09733_ (.A(\instr[6] ),
    .B(\instr[5] ),
    .Y(_04040_));
 sky130_fd_sc_hd__and4b_2 _09734_ (.A_N(_01530_),
    .B(_01854_),
    .C(_04040_),
    .D(\core_state[1] ),
    .X(_04041_));
 sky130_fd_sc_hd__buf_4 _09735_ (.A(_04041_),
    .X(_04042_));
 sky130_fd_sc_hd__or2_4 _09736_ (.A(\core_state[0] ),
    .B(_04042_),
    .X(_04043_));
 sky130_fd_sc_hd__clkbuf_1 _09737_ (.A(_04043_),
    .X(net61));
 sky130_fd_sc_hd__or4bb_1 _09738_ (.A(\instr[3] ),
    .B(\instr[2] ),
    .C_N(\instr[1] ),
    .D_N(\instr[0] ),
    .X(_04044_));
 sky130_fd_sc_hd__buf_4 _09739_ (.A(_04044_),
    .X(_04045_));
 sky130_fd_sc_hd__or4b_4 _09740_ (.A(_01527_),
    .B(\instr[6] ),
    .C(_01530_),
    .D_N(\instr[5] ),
    .X(_04046_));
 sky130_fd_sc_hd__nor2_4 _09741_ (.A(_04045_),
    .B(_04046_),
    .Y(_04047_));
 sky130_fd_sc_hd__buf_4 _09742_ (.A(_04047_),
    .X(_04048_));
 sky130_fd_sc_hd__buf_6 _09743_ (.A(_04048_),
    .X(_04049_));
 sky130_fd_sc_hd__nand2_2 _09744_ (.A(_01642_),
    .B(_01807_),
    .Y(_04050_));
 sky130_fd_sc_hd__or2_1 _09745_ (.A(_01642_),
    .B(_01807_),
    .X(_04051_));
 sky130_fd_sc_hd__and2_2 _09746_ (.A(_04050_),
    .B(_04051_),
    .X(_04052_));
 sky130_fd_sc_hd__or2_1 _09747_ (.A(_01564_),
    .B(_01807_),
    .X(_04053_));
 sky130_fd_sc_hd__and2_1 _09748_ (.A(_01903_),
    .B(_04053_),
    .X(_04054_));
 sky130_fd_sc_hd__a22o_2 _09749_ (.A1(_04049_),
    .A2(_04052_),
    .B1(_04054_),
    .B2(_04042_),
    .X(net37));
 sky130_fd_sc_hd__xor2_4 _09750_ (.A(\B_type_imm[1] ),
    .B(\leorv32_alu.input1[1] ),
    .X(_04055_));
 sky130_fd_sc_hd__xnor2_4 _09751_ (.A(_04050_),
    .B(_04055_),
    .Y(_04056_));
 sky130_fd_sc_hd__buf_6 _09752_ (.A(_04047_),
    .X(_04057_));
 sky130_fd_sc_hd__mux2_1 _09753_ (.A0(\PC[1] ),
    .A1(_04056_),
    .S(_04057_),
    .X(_04058_));
 sky130_fd_sc_hd__clkinv_4 _09754_ (.A(_04041_),
    .Y(_04059_));
 sky130_fd_sc_hd__buf_4 _09755_ (.A(_04059_),
    .X(_04060_));
 sky130_fd_sc_hd__mux2_2 _09756_ (.A0(_04034_),
    .A1(_04058_),
    .S(_04060_),
    .X(_04061_));
 sky130_fd_sc_hd__clkbuf_1 _09757_ (.A(_04061_),
    .X(net48));
 sky130_fd_sc_hd__buf_4 _09758_ (.A(_04060_),
    .X(_04062_));
 sky130_fd_sc_hd__and2_1 _09759_ (.A(\B_type_imm[1] ),
    .B(\leorv32_alu.input1[1] ),
    .X(_04063_));
 sky130_fd_sc_hd__a31oi_4 _09760_ (.A1(\B_type_imm[11] ),
    .A2(\leorv32_alu.input1[0] ),
    .A3(_04055_),
    .B1(_04063_),
    .Y(_04064_));
 sky130_fd_sc_hd__nor2_1 _09761_ (.A(\B_type_imm[2] ),
    .B(_01901_),
    .Y(_04065_));
 sky130_fd_sc_hd__nand2_1 _09762_ (.A(\B_type_imm[2] ),
    .B(_01901_),
    .Y(_04066_));
 sky130_fd_sc_hd__and2b_1 _09763_ (.A_N(_04065_),
    .B(_04066_),
    .X(_04067_));
 sky130_fd_sc_hd__nand2_1 _09764_ (.A(_04064_),
    .B(_04067_),
    .Y(_04068_));
 sky130_fd_sc_hd__o21a_1 _09765_ (.A1(_04064_),
    .A2(_04067_),
    .B1(_04057_),
    .X(_04069_));
 sky130_fd_sc_hd__nor2_1 _09766_ (.A(_01585_),
    .B(_04048_),
    .Y(_04070_));
 sky130_fd_sc_hd__a211o_1 _09767_ (.A1(_04068_),
    .A2(_04069_),
    .B1(_04070_),
    .C1(_04042_),
    .X(_04071_));
 sky130_fd_sc_hd__o21ai_2 _09768_ (.A1(_02246_),
    .A2(_04062_),
    .B1(_04071_),
    .Y(net53));
 sky130_fd_sc_hd__nor2_1 _09769_ (.A(_02315_),
    .B(_01898_),
    .Y(_04072_));
 sky130_fd_sc_hd__nand2_1 _09770_ (.A(_02315_),
    .B(_01898_),
    .Y(_04073_));
 sky130_fd_sc_hd__or2b_1 _09771_ (.A(_04072_),
    .B_N(_04073_),
    .X(_04074_));
 sky130_fd_sc_hd__o21ai_1 _09772_ (.A1(_04064_),
    .A2(_04065_),
    .B1(_04066_),
    .Y(_04075_));
 sky130_fd_sc_hd__xnor2_1 _09773_ (.A(_04074_),
    .B(_04075_),
    .Y(_04076_));
 sky130_fd_sc_hd__mux2_1 _09774_ (.A0(\PC[3] ),
    .A1(_04076_),
    .S(_04057_),
    .X(_04077_));
 sky130_fd_sc_hd__mux2_2 _09775_ (.A0(_02235_),
    .A1(_04077_),
    .S(_04060_),
    .X(_04078_));
 sky130_fd_sc_hd__clkbuf_1 _09776_ (.A(_04078_),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_4 _09777_ (.A(_04057_),
    .X(_04079_));
 sky130_fd_sc_hd__nor2_1 _09778_ (.A(\B_type_imm[4] ),
    .B(_01764_),
    .Y(_04080_));
 sky130_fd_sc_hd__nand2_1 _09779_ (.A(_02313_),
    .B(_01764_),
    .Y(_04081_));
 sky130_fd_sc_hd__or2b_1 _09780_ (.A(_04080_),
    .B_N(_04081_),
    .X(_04082_));
 sky130_fd_sc_hd__o211a_1 _09781_ (.A1(_04064_),
    .A2(_04065_),
    .B1(_04066_),
    .C1(_04073_),
    .X(_04083_));
 sky130_fd_sc_hd__or2_1 _09782_ (.A(_04072_),
    .B(_04083_),
    .X(_04084_));
 sky130_fd_sc_hd__xnor2_1 _09783_ (.A(_04082_),
    .B(_04084_),
    .Y(_04085_));
 sky130_fd_sc_hd__nor2_1 _09784_ (.A(\PC[4] ),
    .B(_04048_),
    .Y(_04086_));
 sky130_fd_sc_hd__a211o_1 _09785_ (.A1(_04079_),
    .A2(_04085_),
    .B1(_04086_),
    .C1(_04042_),
    .X(_04087_));
 sky130_fd_sc_hd__o21ai_2 _09786_ (.A1(_02221_),
    .A2(_04062_),
    .B1(_04087_),
    .Y(net55));
 sky130_fd_sc_hd__o31ai_2 _09787_ (.A1(_04072_),
    .A2(_04080_),
    .A3(_04083_),
    .B1(_04081_),
    .Y(_04088_));
 sky130_fd_sc_hd__xor2_1 _09788_ (.A(_01912_),
    .B(_04088_),
    .X(_04089_));
 sky130_fd_sc_hd__nor2_1 _09789_ (.A(\PC[5] ),
    .B(_04048_),
    .Y(_04090_));
 sky130_fd_sc_hd__a211o_1 _09790_ (.A1(_04079_),
    .A2(_04089_),
    .B1(_04090_),
    .C1(_04042_),
    .X(_04091_));
 sky130_fd_sc_hd__o21ai_1 _09791_ (.A1(_02208_),
    .A2(_04062_),
    .B1(_04091_),
    .Y(net56));
 sky130_fd_sc_hd__a21boi_1 _09792_ (.A1(_01911_),
    .A2(_04088_),
    .B1_N(_01891_),
    .Y(_04092_));
 sky130_fd_sc_hd__xnor2_1 _09793_ (.A(_01915_),
    .B(_04092_),
    .Y(_04093_));
 sky130_fd_sc_hd__nor2_1 _09794_ (.A(_01591_),
    .B(_04048_),
    .Y(_04094_));
 sky130_fd_sc_hd__a211o_1 _09795_ (.A1(_04079_),
    .A2(_04093_),
    .B1(_04094_),
    .C1(_04042_),
    .X(_04095_));
 sky130_fd_sc_hd__o21ai_1 _09796_ (.A1(_02196_),
    .A2(_04062_),
    .B1(_04095_),
    .Y(net57));
 sky130_fd_sc_hd__o21a_1 _09797_ (.A1(_01915_),
    .A2(_04092_),
    .B1(_01889_),
    .X(_04096_));
 sky130_fd_sc_hd__and2_1 _09798_ (.A(_02185_),
    .B(_04096_),
    .X(_04097_));
 sky130_fd_sc_hd__o21ai_1 _09799_ (.A1(_02185_),
    .A2(_04096_),
    .B1(_04079_),
    .Y(_04098_));
 sky130_fd_sc_hd__o221ai_1 _09800_ (.A1(\PC[7] ),
    .A2(_04049_),
    .B1(_04097_),
    .B2(_04098_),
    .C1(_04060_),
    .Y(_04099_));
 sky130_fd_sc_hd__o21ai_1 _09801_ (.A1(_02186_),
    .A2(_04062_),
    .B1(_04099_),
    .Y(net58));
 sky130_fd_sc_hd__o21ai_1 _09802_ (.A1(_01921_),
    .A2(_04096_),
    .B1(_01888_),
    .Y(_04100_));
 sky130_fd_sc_hd__xnor2_1 _09803_ (.A(_01920_),
    .B(_04100_),
    .Y(_04101_));
 sky130_fd_sc_hd__mux2_1 _09804_ (.A0(\PC[8] ),
    .A1(_04101_),
    .S(_04057_),
    .X(_04102_));
 sky130_fd_sc_hd__mux2_1 _09805_ (.A0(_02177_),
    .A1(_04102_),
    .S(_04060_),
    .X(_04103_));
 sky130_fd_sc_hd__clkbuf_1 _09806_ (.A(_04103_),
    .X(net59));
 sky130_fd_sc_hd__and2b_1 _09807_ (.A_N(_01920_),
    .B(_04100_),
    .X(_04104_));
 sky130_fd_sc_hd__nor2_1 _09808_ (.A(_01918_),
    .B(_04104_),
    .Y(_04105_));
 sky130_fd_sc_hd__xnor2_1 _09809_ (.A(_01886_),
    .B(_04105_),
    .Y(_04106_));
 sky130_fd_sc_hd__mux2_1 _09810_ (.A0(\PC[9] ),
    .A1(_04106_),
    .S(_04057_),
    .X(_04107_));
 sky130_fd_sc_hd__mux2_1 _09811_ (.A0(_02155_),
    .A1(_04107_),
    .S(_04060_),
    .X(_04108_));
 sky130_fd_sc_hd__clkbuf_1 _09812_ (.A(_04108_),
    .X(net60));
 sky130_fd_sc_hd__o31a_1 _09813_ (.A1(_01883_),
    .A2(_01918_),
    .A3(_04104_),
    .B1(_01884_),
    .X(_04109_));
 sky130_fd_sc_hd__xor2_1 _09814_ (.A(_01882_),
    .B(_04109_),
    .X(_04110_));
 sky130_fd_sc_hd__mux2_1 _09815_ (.A0(\PC[10] ),
    .A1(_04110_),
    .S(_04057_),
    .X(_04111_));
 sky130_fd_sc_hd__mux2_1 _09816_ (.A0(_02146_),
    .A1(_04111_),
    .S(_04059_),
    .X(_04112_));
 sky130_fd_sc_hd__clkbuf_1 _09817_ (.A(_04112_),
    .X(net38));
 sky130_fd_sc_hd__a21oi_1 _09818_ (.A1(_01882_),
    .A2(_04109_),
    .B1(_01881_),
    .Y(_04113_));
 sky130_fd_sc_hd__xnor2_1 _09819_ (.A(_01876_),
    .B(_04113_),
    .Y(_04114_));
 sky130_fd_sc_hd__mux2_1 _09820_ (.A0(\PC[11] ),
    .A1(_04114_),
    .S(_04079_),
    .X(_04115_));
 sky130_fd_sc_hd__nor2_1 _09821_ (.A(_02134_),
    .B(_04060_),
    .Y(_04116_));
 sky130_fd_sc_hd__a21o_1 _09822_ (.A1(_04062_),
    .A2(_04115_),
    .B1(_04116_),
    .X(net39));
 sky130_fd_sc_hd__a41oi_4 _09823_ (.A1(_01876_),
    .A2(_01882_),
    .A3(_01886_),
    .A4(_04104_),
    .B1(_01926_),
    .Y(_04117_));
 sky130_fd_sc_hd__xnor2_1 _09824_ (.A(_01931_),
    .B(_04117_),
    .Y(_04118_));
 sky130_fd_sc_hd__nor2_1 _09825_ (.A(_01558_),
    .B(_04048_),
    .Y(_04119_));
 sky130_fd_sc_hd__a211o_1 _09826_ (.A1(_04079_),
    .A2(_04118_),
    .B1(_04119_),
    .C1(_04042_),
    .X(_04120_));
 sky130_fd_sc_hd__o21ai_1 _09827_ (.A1(_02122_),
    .A2(_04062_),
    .B1(_04120_),
    .Y(net40));
 sky130_fd_sc_hd__nor2_1 _09828_ (.A(_01931_),
    .B(_04117_),
    .Y(_04121_));
 sky130_fd_sc_hd__or3_1 _09829_ (.A(_01928_),
    .B(_01932_),
    .C(_04121_),
    .X(_04122_));
 sky130_fd_sc_hd__o21ai_1 _09830_ (.A1(_01928_),
    .A2(_04121_),
    .B1(_01932_),
    .Y(_04123_));
 sky130_fd_sc_hd__o21a_1 _09831_ (.A1(_04045_),
    .A2(_04046_),
    .B1(\PC[13] ),
    .X(_04124_));
 sky130_fd_sc_hd__a31o_1 _09832_ (.A1(_04057_),
    .A2(_04122_),
    .A3(_04123_),
    .B1(_04124_),
    .X(_04125_));
 sky130_fd_sc_hd__mux2_1 _09833_ (.A0(_02104_),
    .A1(_04125_),
    .S(_04059_),
    .X(_04126_));
 sky130_fd_sc_hd__clkbuf_1 _09834_ (.A(_04126_),
    .X(net41));
 sky130_fd_sc_hd__a22oi_2 _09835_ (.A1(_01540_),
    .A2(_01873_),
    .B1(_01932_),
    .B2(_04121_),
    .Y(_04127_));
 sky130_fd_sc_hd__xnor2_1 _09836_ (.A(_01936_),
    .B(_04127_),
    .Y(_04128_));
 sky130_fd_sc_hd__nor2_1 _09837_ (.A(\PC[14] ),
    .B(_04048_),
    .Y(_04129_));
 sky130_fd_sc_hd__a211o_1 _09838_ (.A1(_04079_),
    .A2(_04128_),
    .B1(_04129_),
    .C1(_04042_),
    .X(_04130_));
 sky130_fd_sc_hd__o21ai_1 _09839_ (.A1(_02097_),
    .A2(_04062_),
    .B1(_04130_),
    .Y(net42));
 sky130_fd_sc_hd__o21a_1 _09840_ (.A1(_01936_),
    .A2(_04127_),
    .B1(_01934_),
    .X(_04131_));
 sky130_fd_sc_hd__xnor2_1 _09841_ (.A(_01937_),
    .B(_04131_),
    .Y(_04132_));
 sky130_fd_sc_hd__nor2_1 _09842_ (.A(_01615_),
    .B(_04048_),
    .Y(_04133_));
 sky130_fd_sc_hd__a211o_1 _09843_ (.A1(_04079_),
    .A2(_04132_),
    .B1(_04133_),
    .C1(_04042_),
    .X(_04134_));
 sky130_fd_sc_hd__o21ai_1 _09844_ (.A1(_02080_),
    .A2(_04062_),
    .B1(_04134_),
    .Y(net43));
 sky130_fd_sc_hd__nor2_1 _09845_ (.A(_01938_),
    .B(_04117_),
    .Y(_04135_));
 sky130_fd_sc_hd__nor3_1 _09846_ (.A(_01942_),
    .B(_01875_),
    .C(_04135_),
    .Y(_04136_));
 sky130_fd_sc_hd__o21a_1 _09847_ (.A1(_01875_),
    .A2(_04135_),
    .B1(_01942_),
    .X(_04137_));
 sky130_fd_sc_hd__o21ai_1 _09848_ (.A1(_04136_),
    .A2(_04137_),
    .B1(_04049_),
    .Y(_04138_));
 sky130_fd_sc_hd__clkbuf_4 _09849_ (.A(_04057_),
    .X(_04139_));
 sky130_fd_sc_hd__o21a_1 _09850_ (.A1(\PC[16] ),
    .A2(_04139_),
    .B1(_04060_),
    .X(_04140_));
 sky130_fd_sc_hd__a2bb2o_1 _09851_ (.A1_N(_02063_),
    .A2_N(_04062_),
    .B1(_04138_),
    .B2(_04140_),
    .X(net44));
 sky130_fd_sc_hd__or2_1 _09852_ (.A(_01940_),
    .B(_04137_),
    .X(_04141_));
 sky130_fd_sc_hd__xnor2_1 _09853_ (.A(_01944_),
    .B(_04141_),
    .Y(_04142_));
 sky130_fd_sc_hd__nor2_1 _09854_ (.A(\PC[17] ),
    .B(_04048_),
    .Y(_04143_));
 sky130_fd_sc_hd__a211o_1 _09855_ (.A1(_04079_),
    .A2(_04142_),
    .B1(_04143_),
    .C1(_04042_),
    .X(_04144_));
 sky130_fd_sc_hd__o21ai_1 _09856_ (.A1(_02049_),
    .A2(_04060_),
    .B1(_04144_),
    .Y(net45));
 sky130_fd_sc_hd__nand2_1 _09857_ (.A(_01944_),
    .B(_04137_),
    .Y(_04145_));
 sky130_fd_sc_hd__and3_1 _09858_ (.A(_01946_),
    .B(_02023_),
    .C(_04145_),
    .X(_04146_));
 sky130_fd_sc_hd__a21oi_1 _09859_ (.A1(_02023_),
    .A2(_04145_),
    .B1(_01946_),
    .Y(_04147_));
 sky130_fd_sc_hd__o21ai_1 _09860_ (.A1(_04045_),
    .A2(_04046_),
    .B1(\PC[18] ),
    .Y(_04148_));
 sky130_fd_sc_hd__o41ai_1 _09861_ (.A1(_04045_),
    .A2(_04046_),
    .A3(_04146_),
    .A4(_04147_),
    .B1(_04148_),
    .Y(_04149_));
 sky130_fd_sc_hd__mux2_1 _09862_ (.A0(_02032_),
    .A1(_04149_),
    .S(_04059_),
    .X(_04150_));
 sky130_fd_sc_hd__clkbuf_1 _09863_ (.A(_04150_),
    .X(net46));
 sky130_fd_sc_hd__a21oi_1 _09864_ (.A1(_01540_),
    .A2(_01867_),
    .B1(_04147_),
    .Y(_04151_));
 sky130_fd_sc_hd__xnor2_1 _09865_ (.A(_01947_),
    .B(_04151_),
    .Y(_04152_));
 sky130_fd_sc_hd__mux2_1 _09866_ (.A0(\PC[19] ),
    .A1(_04152_),
    .S(_04047_),
    .X(_04153_));
 sky130_fd_sc_hd__mux2_1 _09867_ (.A0(_02026_),
    .A1(_04153_),
    .S(_04059_),
    .X(_04154_));
 sky130_fd_sc_hd__clkbuf_1 _09868_ (.A(_04154_),
    .X(net47));
 sky130_fd_sc_hd__o2bb2a_1 _09869_ (.A1_N(_01538_),
    .A2_N(_01869_),
    .B1(_01948_),
    .B2(_04145_),
    .X(_04155_));
 sky130_fd_sc_hd__xnor2_1 _09870_ (.A(_01866_),
    .B(_04155_),
    .Y(_04156_));
 sky130_fd_sc_hd__nor2_1 _09871_ (.A(_01546_),
    .B(_04048_),
    .Y(_04157_));
 sky130_fd_sc_hd__a211o_1 _09872_ (.A1(_04079_),
    .A2(_04156_),
    .B1(_04157_),
    .C1(_04041_),
    .X(_04158_));
 sky130_fd_sc_hd__o21ai_1 _09873_ (.A1(_02011_),
    .A2(_04060_),
    .B1(_04158_),
    .Y(net49));
 sky130_fd_sc_hd__or2_1 _09874_ (.A(_01866_),
    .B(_04155_),
    .X(_04159_));
 sky130_fd_sc_hd__nand2_1 _09875_ (.A(_01864_),
    .B(_04159_),
    .Y(_04160_));
 sky130_fd_sc_hd__xnor2_1 _09876_ (.A(_01951_),
    .B(_04160_),
    .Y(_04161_));
 sky130_fd_sc_hd__mux2_1 _09877_ (.A0(\PC[21] ),
    .A1(_04161_),
    .S(_04047_),
    .X(_04162_));
 sky130_fd_sc_hd__mux2_1 _09878_ (.A0(_01988_),
    .A1(_04162_),
    .S(_04059_),
    .X(_04163_));
 sky130_fd_sc_hd__clkbuf_1 _09879_ (.A(_04163_),
    .X(net50));
 sky130_fd_sc_hd__o2bb2a_1 _09880_ (.A1_N(_01539_),
    .A2_N(_01863_),
    .B1(_04159_),
    .B2(_01951_),
    .X(_04164_));
 sky130_fd_sc_hd__xnor2_1 _09881_ (.A(_01963_),
    .B(_04164_),
    .Y(_04165_));
 sky130_fd_sc_hd__mux2_1 _09882_ (.A0(\PC[22] ),
    .A1(_04165_),
    .S(_04047_),
    .X(_04166_));
 sky130_fd_sc_hd__mux2_1 _09883_ (.A0(_01964_),
    .A1(_04166_),
    .S(_04059_),
    .X(_04167_));
 sky130_fd_sc_hd__clkbuf_1 _09884_ (.A(_04167_),
    .X(net51));
 sky130_fd_sc_hd__o21ai_1 _09885_ (.A1(_01862_),
    .A2(_04164_),
    .B1(_01953_),
    .Y(_04168_));
 sky130_fd_sc_hd__xnor2_1 _09886_ (.A(_01955_),
    .B(_04168_),
    .Y(_04169_));
 sky130_fd_sc_hd__mux2_1 _09887_ (.A0(\PC[23] ),
    .A1(_04169_),
    .S(_04047_),
    .X(_04170_));
 sky130_fd_sc_hd__mux2_1 _09888_ (.A0(_01956_),
    .A1(_04170_),
    .S(_04059_),
    .X(_04171_));
 sky130_fd_sc_hd__clkbuf_1 _09889_ (.A(_04171_),
    .X(net52));
 sky130_fd_sc_hd__or2_1 _09890_ (.A(_01826_),
    .B(_01979_),
    .X(_04172_));
 sky130_fd_sc_hd__buf_4 _09891_ (.A(_04172_),
    .X(_04173_));
 sky130_fd_sc_hd__o21a_2 _09892_ (.A1(_04052_),
    .A2(_04056_),
    .B1(_04173_),
    .X(_04174_));
 sky130_fd_sc_hd__a2111o_4 _09893_ (.A1(_01689_),
    .A2(_01826_),
    .B1(_04045_),
    .C1(_04046_),
    .D1(_02308_),
    .X(_04175_));
 sky130_fd_sc_hd__nor2_8 _09894_ (.A(_04174_),
    .B(_04175_),
    .Y(net94));
 sky130_fd_sc_hd__a21oi_4 _09895_ (.A1(_01832_),
    .A2(_04173_),
    .B1(_04174_),
    .Y(_04176_));
 sky130_fd_sc_hd__buf_4 _09896_ (.A(_01824_),
    .X(_04177_));
 sky130_fd_sc_hd__clkbuf_4 _09897_ (.A(_04177_),
    .X(_04178_));
 sky130_fd_sc_hd__and3b_1 _09898_ (.A_N(_04055_),
    .B(_04052_),
    .C(_04178_),
    .X(_04179_));
 sky130_fd_sc_hd__clkbuf_4 _09899_ (.A(_04179_),
    .X(_04180_));
 sky130_fd_sc_hd__o21a_1 _09900_ (.A1(_04176_),
    .A2(_04180_),
    .B1(_04049_),
    .X(net95));
 sky130_fd_sc_hd__or2b_2 _09901_ (.A(_04052_),
    .B_N(_04056_),
    .X(_04181_));
 sky130_fd_sc_hd__a21oi_4 _09902_ (.A1(_04173_),
    .A2(_04181_),
    .B1(_04175_),
    .Y(net96));
 sky130_fd_sc_hd__nor2_2 _09903_ (.A(_01826_),
    .B(_01979_),
    .Y(_04182_));
 sky130_fd_sc_hd__clkbuf_4 _09904_ (.A(_04182_),
    .X(_04183_));
 sky130_fd_sc_hd__buf_2 _09905_ (.A(_04183_),
    .X(_04184_));
 sky130_fd_sc_hd__nor2_2 _09906_ (.A(_01832_),
    .B(_04181_),
    .Y(_04185_));
 sky130_fd_sc_hd__and3_1 _09907_ (.A(_04178_),
    .B(_04052_),
    .C(_04055_),
    .X(_04186_));
 sky130_fd_sc_hd__clkbuf_2 _09908_ (.A(_04186_),
    .X(_04187_));
 sky130_fd_sc_hd__o31a_2 _09909_ (.A1(_04184_),
    .A2(_04185_),
    .A3(_04187_),
    .B1(_04049_),
    .X(net97));
 sky130_fd_sc_hd__and2_1 _09910_ (.A(\rs2_content[0] ),
    .B(net94),
    .X(_04188_));
 sky130_fd_sc_hd__clkbuf_1 _09911_ (.A(_04188_),
    .X(net62));
 sky130_fd_sc_hd__and2_1 _09912_ (.A(\rs2_content[1] ),
    .B(net94),
    .X(_04189_));
 sky130_fd_sc_hd__clkbuf_1 _09913_ (.A(_04189_),
    .X(net73));
 sky130_fd_sc_hd__and2_1 _09914_ (.A(_01772_),
    .B(net94),
    .X(_04190_));
 sky130_fd_sc_hd__clkbuf_1 _09915_ (.A(_04190_),
    .X(net84));
 sky130_fd_sc_hd__and2_1 _09916_ (.A(_01770_),
    .B(net94),
    .X(_04191_));
 sky130_fd_sc_hd__clkbuf_1 _09917_ (.A(_04191_),
    .X(net87));
 sky130_fd_sc_hd__and2_1 _09918_ (.A(\rs2_content[4] ),
    .B(net94),
    .X(_04192_));
 sky130_fd_sc_hd__clkbuf_1 _09919_ (.A(_04192_),
    .X(net88));
 sky130_fd_sc_hd__and2_1 _09920_ (.A(\rs2_content[5] ),
    .B(net94),
    .X(_04193_));
 sky130_fd_sc_hd__clkbuf_1 _09921_ (.A(_04193_),
    .X(net89));
 sky130_fd_sc_hd__and2_1 _09922_ (.A(\rs2_content[6] ),
    .B(net94),
    .X(_04194_));
 sky130_fd_sc_hd__clkbuf_1 _09923_ (.A(_04194_),
    .X(net90));
 sky130_fd_sc_hd__and2_1 _09924_ (.A(\rs2_content[7] ),
    .B(net94),
    .X(_04195_));
 sky130_fd_sc_hd__clkbuf_1 _09925_ (.A(_04195_),
    .X(net91));
 sky130_fd_sc_hd__a22o_1 _09926_ (.A1(\rs2_content[8] ),
    .A2(_04176_),
    .B1(_04180_),
    .B2(\rs2_content[0] ),
    .X(_04196_));
 sky130_fd_sc_hd__and2_1 _09927_ (.A(_04049_),
    .B(_04196_),
    .X(_04197_));
 sky130_fd_sc_hd__clkbuf_1 _09928_ (.A(_04197_),
    .X(net92));
 sky130_fd_sc_hd__a22o_1 _09929_ (.A1(\rs2_content[9] ),
    .A2(_04176_),
    .B1(_04180_),
    .B2(\rs2_content[1] ),
    .X(_04198_));
 sky130_fd_sc_hd__and2_1 _09930_ (.A(_04049_),
    .B(_04198_),
    .X(_04199_));
 sky130_fd_sc_hd__clkbuf_1 _09931_ (.A(_04199_),
    .X(net93));
 sky130_fd_sc_hd__a22o_1 _09932_ (.A1(\rs2_content[10] ),
    .A2(_04176_),
    .B1(_04180_),
    .B2(_01772_),
    .X(_04200_));
 sky130_fd_sc_hd__and2_1 _09933_ (.A(_04049_),
    .B(_04200_),
    .X(_04201_));
 sky130_fd_sc_hd__clkbuf_1 _09934_ (.A(_04201_),
    .X(net63));
 sky130_fd_sc_hd__a22o_1 _09935_ (.A1(\rs2_content[11] ),
    .A2(_04176_),
    .B1(_04180_),
    .B2(_01770_),
    .X(_04202_));
 sky130_fd_sc_hd__and2_1 _09936_ (.A(_04049_),
    .B(_04202_),
    .X(_04203_));
 sky130_fd_sc_hd__clkbuf_1 _09937_ (.A(_04203_),
    .X(net64));
 sky130_fd_sc_hd__buf_2 _09938_ (.A(_04057_),
    .X(_04204_));
 sky130_fd_sc_hd__a22o_1 _09939_ (.A1(\rs2_content[12] ),
    .A2(_04176_),
    .B1(_04180_),
    .B2(\rs2_content[4] ),
    .X(_04205_));
 sky130_fd_sc_hd__and2_1 _09940_ (.A(_04204_),
    .B(_04205_),
    .X(_04206_));
 sky130_fd_sc_hd__clkbuf_1 _09941_ (.A(_04206_),
    .X(net65));
 sky130_fd_sc_hd__a22o_1 _09942_ (.A1(\rs2_content[13] ),
    .A2(_04176_),
    .B1(_04180_),
    .B2(\rs2_content[5] ),
    .X(_04207_));
 sky130_fd_sc_hd__and2_1 _09943_ (.A(_04204_),
    .B(_04207_),
    .X(_04208_));
 sky130_fd_sc_hd__clkbuf_1 _09944_ (.A(_04208_),
    .X(net66));
 sky130_fd_sc_hd__a22o_1 _09945_ (.A1(\rs2_content[14] ),
    .A2(_04176_),
    .B1(_04180_),
    .B2(\rs2_content[6] ),
    .X(_04209_));
 sky130_fd_sc_hd__and2_1 _09946_ (.A(_04204_),
    .B(_04209_),
    .X(_04210_));
 sky130_fd_sc_hd__clkbuf_1 _09947_ (.A(_04210_),
    .X(net67));
 sky130_fd_sc_hd__a22o_1 _09948_ (.A1(\rs2_content[15] ),
    .A2(_04176_),
    .B1(_04180_),
    .B2(\rs2_content[7] ),
    .X(_04211_));
 sky130_fd_sc_hd__and2_1 _09949_ (.A(_04204_),
    .B(_04211_),
    .X(_04212_));
 sky130_fd_sc_hd__clkbuf_1 _09950_ (.A(_04212_),
    .X(net68));
 sky130_fd_sc_hd__nor3_4 _09951_ (.A(_02308_),
    .B(_01689_),
    .C(_04181_),
    .Y(_04213_));
 sky130_fd_sc_hd__a22o_1 _09952_ (.A1(\rs2_content[16] ),
    .A2(_04184_),
    .B1(_04213_),
    .B2(\rs2_content[0] ),
    .X(_04214_));
 sky130_fd_sc_hd__and2_1 _09953_ (.A(_04204_),
    .B(_04214_),
    .X(_04215_));
 sky130_fd_sc_hd__clkbuf_1 _09954_ (.A(_04215_),
    .X(net69));
 sky130_fd_sc_hd__a22o_1 _09955_ (.A1(\rs2_content[17] ),
    .A2(_04184_),
    .B1(_04213_),
    .B2(\rs2_content[1] ),
    .X(_04216_));
 sky130_fd_sc_hd__and2_1 _09956_ (.A(_04204_),
    .B(_04216_),
    .X(_04217_));
 sky130_fd_sc_hd__clkbuf_1 _09957_ (.A(_04217_),
    .X(net70));
 sky130_fd_sc_hd__a22o_1 _09958_ (.A1(\rs2_content[18] ),
    .A2(_04184_),
    .B1(_04213_),
    .B2(_01772_),
    .X(_04218_));
 sky130_fd_sc_hd__and2_1 _09959_ (.A(_04204_),
    .B(_04218_),
    .X(_04219_));
 sky130_fd_sc_hd__clkbuf_1 _09960_ (.A(_04219_),
    .X(net71));
 sky130_fd_sc_hd__a22o_1 _09961_ (.A1(\rs2_content[19] ),
    .A2(_04184_),
    .B1(_04213_),
    .B2(_01770_),
    .X(_04220_));
 sky130_fd_sc_hd__and2_1 _09962_ (.A(_04204_),
    .B(_04220_),
    .X(_04221_));
 sky130_fd_sc_hd__clkbuf_1 _09963_ (.A(_04221_),
    .X(net72));
 sky130_fd_sc_hd__a22o_1 _09964_ (.A1(\rs2_content[20] ),
    .A2(_04184_),
    .B1(_04213_),
    .B2(\rs2_content[4] ),
    .X(_04222_));
 sky130_fd_sc_hd__and2_1 _09965_ (.A(_04204_),
    .B(_04222_),
    .X(_04223_));
 sky130_fd_sc_hd__clkbuf_1 _09966_ (.A(_04223_),
    .X(net74));
 sky130_fd_sc_hd__a22o_1 _09967_ (.A1(\rs2_content[21] ),
    .A2(_04184_),
    .B1(_04213_),
    .B2(\rs2_content[5] ),
    .X(_04224_));
 sky130_fd_sc_hd__and2_1 _09968_ (.A(_04204_),
    .B(_04224_),
    .X(_04225_));
 sky130_fd_sc_hd__clkbuf_1 _09969_ (.A(_04225_),
    .X(net75));
 sky130_fd_sc_hd__a22o_1 _09970_ (.A1(\rs2_content[22] ),
    .A2(_04184_),
    .B1(_04213_),
    .B2(\rs2_content[6] ),
    .X(_04226_));
 sky130_fd_sc_hd__and2_1 _09971_ (.A(_04139_),
    .B(_04226_),
    .X(_04227_));
 sky130_fd_sc_hd__clkbuf_1 _09972_ (.A(_04227_),
    .X(net76));
 sky130_fd_sc_hd__a22o_1 _09973_ (.A1(\rs2_content[23] ),
    .A2(_04184_),
    .B1(_04213_),
    .B2(\rs2_content[7] ),
    .X(_04228_));
 sky130_fd_sc_hd__and2_1 _09974_ (.A(_04139_),
    .B(_04228_),
    .X(_04229_));
 sky130_fd_sc_hd__clkbuf_1 _09975_ (.A(_04229_),
    .X(net77));
 sky130_fd_sc_hd__a22o_1 _09976_ (.A1(\rs2_content[24] ),
    .A2(_04184_),
    .B1(_04187_),
    .B2(\rs2_content[0] ),
    .X(_04230_));
 sky130_fd_sc_hd__a21o_1 _09977_ (.A1(\rs2_content[8] ),
    .A2(_04185_),
    .B1(_04230_),
    .X(_04231_));
 sky130_fd_sc_hd__and2_1 _09978_ (.A(_04139_),
    .B(_04231_),
    .X(_04232_));
 sky130_fd_sc_hd__clkbuf_1 _09979_ (.A(_04232_),
    .X(net78));
 sky130_fd_sc_hd__a22o_1 _09980_ (.A1(\rs2_content[25] ),
    .A2(_04183_),
    .B1(_04187_),
    .B2(\rs2_content[1] ),
    .X(_04233_));
 sky130_fd_sc_hd__a21o_1 _09981_ (.A1(\rs2_content[9] ),
    .A2(_04185_),
    .B1(_04233_),
    .X(_04234_));
 sky130_fd_sc_hd__and2_1 _09982_ (.A(_04139_),
    .B(_04234_),
    .X(_04235_));
 sky130_fd_sc_hd__clkbuf_1 _09983_ (.A(_04235_),
    .X(net79));
 sky130_fd_sc_hd__nor2_1 _09984_ (.A(_01707_),
    .B(_04173_),
    .Y(_04236_));
 sky130_fd_sc_hd__a22o_1 _09985_ (.A1(\rs2_content[10] ),
    .A2(_04185_),
    .B1(_04187_),
    .B2(_01772_),
    .X(_04237_));
 sky130_fd_sc_hd__o21a_1 _09986_ (.A1(_04236_),
    .A2(_04237_),
    .B1(_04049_),
    .X(net80));
 sky130_fd_sc_hd__a22o_1 _09987_ (.A1(\rs2_content[27] ),
    .A2(_04183_),
    .B1(_04187_),
    .B2(_01770_),
    .X(_04238_));
 sky130_fd_sc_hd__a21o_1 _09988_ (.A1(\rs2_content[11] ),
    .A2(_04185_),
    .B1(_04238_),
    .X(_04239_));
 sky130_fd_sc_hd__and2_1 _09989_ (.A(_04139_),
    .B(_04239_),
    .X(_04240_));
 sky130_fd_sc_hd__clkbuf_1 _09990_ (.A(_04240_),
    .X(net81));
 sky130_fd_sc_hd__a22o_1 _09991_ (.A1(\rs2_content[28] ),
    .A2(_04183_),
    .B1(_04187_),
    .B2(\rs2_content[4] ),
    .X(_04241_));
 sky130_fd_sc_hd__a21o_1 _09992_ (.A1(\rs2_content[12] ),
    .A2(_04185_),
    .B1(_04241_),
    .X(_04242_));
 sky130_fd_sc_hd__and2_1 _09993_ (.A(_04139_),
    .B(_04242_),
    .X(_04243_));
 sky130_fd_sc_hd__clkbuf_1 _09994_ (.A(_04243_),
    .X(net82));
 sky130_fd_sc_hd__a22o_1 _09995_ (.A1(\rs2_content[29] ),
    .A2(_04183_),
    .B1(_04187_),
    .B2(\rs2_content[5] ),
    .X(_04244_));
 sky130_fd_sc_hd__a21o_1 _09996_ (.A1(\rs2_content[13] ),
    .A2(_04185_),
    .B1(_04244_),
    .X(_04245_));
 sky130_fd_sc_hd__and2_1 _09997_ (.A(_04139_),
    .B(_04245_),
    .X(_04246_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _09998_ (.A(_04246_),
    .X(net83));
 sky130_fd_sc_hd__a22o_1 _09999_ (.A1(\rs2_content[30] ),
    .A2(_04183_),
    .B1(_04187_),
    .B2(\rs2_content[6] ),
    .X(_04247_));
 sky130_fd_sc_hd__a21o_1 _10000_ (.A1(\rs2_content[14] ),
    .A2(_04185_),
    .B1(_04247_),
    .X(_04248_));
 sky130_fd_sc_hd__and2_1 _10001_ (.A(_04139_),
    .B(_04248_),
    .X(_04249_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _10002_ (.A(_04249_),
    .X(net85));
 sky130_fd_sc_hd__a22o_1 _10003_ (.A1(\rs2_content[31] ),
    .A2(_04183_),
    .B1(_04187_),
    .B2(\rs2_content[7] ),
    .X(_04250_));
 sky130_fd_sc_hd__a21o_1 _10004_ (.A1(\rs2_content[15] ),
    .A2(_04185_),
    .B1(_04250_),
    .X(_04251_));
 sky130_fd_sc_hd__and2_1 _10005_ (.A(_04139_),
    .B(_04251_),
    .X(_04252_));
 sky130_fd_sc_hd__clkbuf_1 _10006_ (.A(_04252_),
    .X(net86));
 sky130_fd_sc_hd__clkinv_2 _10007_ (.A(\cycles[0] ),
    .Y(_00004_));
 sky130_fd_sc_hd__xor2_1 _10008_ (.A(\cycles[0] ),
    .B(\cycles[1] ),
    .X(_00015_));
 sky130_fd_sc_hd__and3_1 _10009_ (.A(\cycles[0] ),
    .B(\cycles[1] ),
    .C(\cycles[2] ),
    .X(_04253_));
 sky130_fd_sc_hd__a21oi_1 _10010_ (.A1(\cycles[0] ),
    .A2(\cycles[1] ),
    .B1(\cycles[2] ),
    .Y(_04254_));
 sky130_fd_sc_hd__nor2_1 _10011_ (.A(_04253_),
    .B(_04254_),
    .Y(_00026_));
 sky130_fd_sc_hd__and4_1 _10012_ (.A(\cycles[0] ),
    .B(\cycles[1] ),
    .C(\cycles[2] ),
    .D(\cycles[3] ),
    .X(_04255_));
 sky130_fd_sc_hd__nor2_1 _10013_ (.A(\cycles[3] ),
    .B(_04253_),
    .Y(_04256_));
 sky130_fd_sc_hd__nor2_1 _10014_ (.A(_04255_),
    .B(_04256_),
    .Y(_00037_));
 sky130_fd_sc_hd__nand2_1 _10015_ (.A(\cycles[4] ),
    .B(_04255_),
    .Y(_04257_));
 sky130_fd_sc_hd__or2_1 _10016_ (.A(\cycles[4] ),
    .B(_04255_),
    .X(_04258_));
 sky130_fd_sc_hd__and2_1 _10017_ (.A(_04257_),
    .B(_04258_),
    .X(_04259_));
 sky130_fd_sc_hd__clkbuf_1 _10018_ (.A(_04259_),
    .X(_00048_));
 sky130_fd_sc_hd__xnor2_1 _10019_ (.A(\cycles[5] ),
    .B(_04257_),
    .Y(_00059_));
 sky130_fd_sc_hd__and4_1 _10020_ (.A(\cycles[4] ),
    .B(\cycles[5] ),
    .C(\cycles[6] ),
    .D(_04255_),
    .X(_04260_));
 sky130_fd_sc_hd__a31o_1 _10021_ (.A1(\cycles[4] ),
    .A2(\cycles[5] ),
    .A3(_04255_),
    .B1(\cycles[6] ),
    .X(_04261_));
 sky130_fd_sc_hd__and2b_1 _10022_ (.A_N(_04260_),
    .B(_04261_),
    .X(_04262_));
 sky130_fd_sc_hd__clkbuf_1 _10023_ (.A(_04262_),
    .X(_00064_));
 sky130_fd_sc_hd__nand2_1 _10024_ (.A(\cycles[7] ),
    .B(_04260_),
    .Y(_04263_));
 sky130_fd_sc_hd__or2_1 _10025_ (.A(\cycles[7] ),
    .B(_04260_),
    .X(_04264_));
 sky130_fd_sc_hd__and2_1 _10026_ (.A(_04263_),
    .B(_04264_),
    .X(_04265_));
 sky130_fd_sc_hd__clkbuf_1 _10027_ (.A(_04265_),
    .X(_00065_));
 sky130_fd_sc_hd__xnor2_1 _10028_ (.A(\cycles[8] ),
    .B(_04263_),
    .Y(_00066_));
 sky130_fd_sc_hd__a31oi_1 _10029_ (.A1(\cycles[7] ),
    .A2(\cycles[8] ),
    .A3(_04260_),
    .B1(\cycles[9] ),
    .Y(_04266_));
 sky130_fd_sc_hd__and4_1 _10030_ (.A(\cycles[7] ),
    .B(\cycles[8] ),
    .C(\cycles[9] ),
    .D(_04260_),
    .X(_04267_));
 sky130_fd_sc_hd__nor2_1 _10031_ (.A(_04266_),
    .B(_04267_),
    .Y(_00067_));
 sky130_fd_sc_hd__xor2_1 _10032_ (.A(\cycles[10] ),
    .B(_04267_),
    .X(_00005_));
 sky130_fd_sc_hd__a21oi_1 _10033_ (.A1(\cycles[10] ),
    .A2(_04267_),
    .B1(\cycles[11] ),
    .Y(_04268_));
 sky130_fd_sc_hd__and3_1 _10034_ (.A(\cycles[10] ),
    .B(\cycles[11] ),
    .C(_04267_),
    .X(_04269_));
 sky130_fd_sc_hd__nor2_1 _10035_ (.A(_04268_),
    .B(_04269_),
    .Y(_00006_));
 sky130_fd_sc_hd__nor2_1 _10036_ (.A(\cycles[12] ),
    .B(_04269_),
    .Y(_04270_));
 sky130_fd_sc_hd__and4_1 _10037_ (.A(\cycles[7] ),
    .B(\cycles[8] ),
    .C(\cycles[9] ),
    .D(_04260_),
    .X(_04271_));
 sky130_fd_sc_hd__and4_1 _10038_ (.A(\cycles[10] ),
    .B(\cycles[11] ),
    .C(\cycles[12] ),
    .D(_04271_),
    .X(_04272_));
 sky130_fd_sc_hd__nor2_1 _10039_ (.A(_04270_),
    .B(_04272_),
    .Y(_00007_));
 sky130_fd_sc_hd__nor2_1 _10040_ (.A(\cycles[13] ),
    .B(_04272_),
    .Y(_04273_));
 sky130_fd_sc_hd__and3_1 _10041_ (.A(\cycles[12] ),
    .B(\cycles[13] ),
    .C(_04269_),
    .X(_04274_));
 sky130_fd_sc_hd__nor2_1 _10042_ (.A(_04273_),
    .B(_04274_),
    .Y(_00008_));
 sky130_fd_sc_hd__xor2_1 _10043_ (.A(\cycles[14] ),
    .B(_04274_),
    .X(_00009_));
 sky130_fd_sc_hd__a21oi_1 _10044_ (.A1(\cycles[14] ),
    .A2(_04274_),
    .B1(\cycles[15] ),
    .Y(_04275_));
 sky130_fd_sc_hd__and3_1 _10045_ (.A(\cycles[14] ),
    .B(\cycles[15] ),
    .C(_04274_),
    .X(_04276_));
 sky130_fd_sc_hd__nor2_1 _10046_ (.A(_04275_),
    .B(_04276_),
    .Y(_00010_));
 sky130_fd_sc_hd__and4_1 _10047_ (.A(\cycles[13] ),
    .B(\cycles[14] ),
    .C(\cycles[15] ),
    .D(_04272_),
    .X(_04277_));
 sky130_fd_sc_hd__xor2_1 _10048_ (.A(\cycles[16] ),
    .B(_04277_),
    .X(_00011_));
 sky130_fd_sc_hd__a21oi_1 _10049_ (.A1(\cycles[16] ),
    .A2(_04277_),
    .B1(\cycles[17] ),
    .Y(_04278_));
 sky130_fd_sc_hd__and3_1 _10050_ (.A(\cycles[16] ),
    .B(\cycles[17] ),
    .C(_04276_),
    .X(_04279_));
 sky130_fd_sc_hd__nor2_1 _10051_ (.A(_04278_),
    .B(_04279_),
    .Y(_00012_));
 sky130_fd_sc_hd__nor2_1 _10052_ (.A(\cycles[18] ),
    .B(_04279_),
    .Y(_04280_));
 sky130_fd_sc_hd__and4_1 _10053_ (.A(\cycles[16] ),
    .B(\cycles[17] ),
    .C(\cycles[18] ),
    .D(_04277_),
    .X(_04281_));
 sky130_fd_sc_hd__nor2_1 _10054_ (.A(_04280_),
    .B(_04281_),
    .Y(_00013_));
 sky130_fd_sc_hd__nor2_1 _10055_ (.A(\cycles[19] ),
    .B(_04281_),
    .Y(_04282_));
 sky130_fd_sc_hd__and4_1 _10056_ (.A(\cycles[16] ),
    .B(\cycles[17] ),
    .C(\cycles[18] ),
    .D(\cycles[19] ),
    .X(_04283_));
 sky130_fd_sc_hd__and4_1 _10057_ (.A(\cycles[14] ),
    .B(\cycles[15] ),
    .C(_04274_),
    .D(_04283_),
    .X(_04284_));
 sky130_fd_sc_hd__nor2_1 _10058_ (.A(_04282_),
    .B(_04284_),
    .Y(_00014_));
 sky130_fd_sc_hd__nor2_1 _10059_ (.A(\cycles[20] ),
    .B(_04284_),
    .Y(_04285_));
 sky130_fd_sc_hd__and3_1 _10060_ (.A(\cycles[19] ),
    .B(\cycles[20] ),
    .C(_04281_),
    .X(_04286_));
 sky130_fd_sc_hd__nor2_1 _10061_ (.A(_04285_),
    .B(_04286_),
    .Y(_00016_));
 sky130_fd_sc_hd__nor2_1 _10062_ (.A(\cycles[21] ),
    .B(_04286_),
    .Y(_04287_));
 sky130_fd_sc_hd__and2_1 _10063_ (.A(\cycles[20] ),
    .B(\cycles[21] ),
    .X(_04288_));
 sky130_fd_sc_hd__and2_1 _10064_ (.A(_04284_),
    .B(_04288_),
    .X(_04289_));
 sky130_fd_sc_hd__nor2_1 _10065_ (.A(_04287_),
    .B(_04289_),
    .Y(_00017_));
 sky130_fd_sc_hd__nor2_1 _10066_ (.A(\cycles[22] ),
    .B(_04289_),
    .Y(_04290_));
 sky130_fd_sc_hd__and3_1 _10067_ (.A(\cycles[21] ),
    .B(\cycles[22] ),
    .C(_04286_),
    .X(_04291_));
 sky130_fd_sc_hd__nor2_1 _10068_ (.A(_04290_),
    .B(_04291_),
    .Y(_00018_));
 sky130_fd_sc_hd__nor2_1 _10069_ (.A(\cycles[23] ),
    .B(_04291_),
    .Y(_04292_));
 sky130_fd_sc_hd__and2_1 _10070_ (.A(\cycles[22] ),
    .B(\cycles[23] ),
    .X(_04293_));
 sky130_fd_sc_hd__and3_1 _10071_ (.A(_04284_),
    .B(_04288_),
    .C(_04293_),
    .X(_04294_));
 sky130_fd_sc_hd__nor2_1 _10072_ (.A(_04292_),
    .B(_04294_),
    .Y(_00019_));
 sky130_fd_sc_hd__nor2_1 _10073_ (.A(\cycles[24] ),
    .B(_04294_),
    .Y(_04295_));
 sky130_fd_sc_hd__nand2_1 _10074_ (.A(\cycles[24] ),
    .B(_04294_),
    .Y(_04296_));
 sky130_fd_sc_hd__and2b_1 _10075_ (.A_N(_04295_),
    .B(_04296_),
    .X(_04297_));
 sky130_fd_sc_hd__clkbuf_1 _10076_ (.A(_04297_),
    .X(_00020_));
 sky130_fd_sc_hd__inv_2 _10077_ (.A(\cycles[25] ),
    .Y(_04298_));
 sky130_fd_sc_hd__and2_1 _10078_ (.A(\cycles[24] ),
    .B(\cycles[25] ),
    .X(_04299_));
 sky130_fd_sc_hd__and4_1 _10079_ (.A(_04284_),
    .B(_04288_),
    .C(_04293_),
    .D(_04299_),
    .X(_04300_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _10080_ (.A(_04300_),
    .X(_04301_));
 sky130_fd_sc_hd__a21oi_1 _10081_ (.A1(_04298_),
    .A2(_04296_),
    .B1(_04301_),
    .Y(_00021_));
 sky130_fd_sc_hd__xor2_1 _10082_ (.A(\cycles[26] ),
    .B(_04301_),
    .X(_00022_));
 sky130_fd_sc_hd__a21oi_1 _10083_ (.A1(\cycles[26] ),
    .A2(_04301_),
    .B1(\cycles[27] ),
    .Y(_04302_));
 sky130_fd_sc_hd__and3_1 _10084_ (.A(\cycles[26] ),
    .B(\cycles[27] ),
    .C(_04301_),
    .X(_04303_));
 sky130_fd_sc_hd__nor2_1 _10085_ (.A(_04302_),
    .B(_04303_),
    .Y(_00023_));
 sky130_fd_sc_hd__xor2_1 _10086_ (.A(\cycles[28] ),
    .B(_04303_),
    .X(_00024_));
 sky130_fd_sc_hd__and4_1 _10087_ (.A(\cycles[23] ),
    .B(\cycles[24] ),
    .C(\cycles[25] ),
    .D(_04291_),
    .X(_04304_));
 sky130_fd_sc_hd__and4_1 _10088_ (.A(\cycles[26] ),
    .B(\cycles[27] ),
    .C(\cycles[28] ),
    .D(_04304_),
    .X(_04305_));
 sky130_fd_sc_hd__xor2_1 _10089_ (.A(\cycles[29] ),
    .B(_04305_),
    .X(_00025_));
 sky130_fd_sc_hd__and2_1 _10090_ (.A(\cycles[28] ),
    .B(\cycles[29] ),
    .X(_04306_));
 sky130_fd_sc_hd__and4_1 _10091_ (.A(\cycles[26] ),
    .B(\cycles[27] ),
    .C(_04301_),
    .D(_04306_),
    .X(_04307_));
 sky130_fd_sc_hd__xor2_1 _10092_ (.A(\cycles[30] ),
    .B(_04307_),
    .X(_00027_));
 sky130_fd_sc_hd__a21oi_1 _10093_ (.A1(\cycles[30] ),
    .A2(_04307_),
    .B1(\cycles[31] ),
    .Y(_04308_));
 sky130_fd_sc_hd__and4_1 _10094_ (.A(\cycles[29] ),
    .B(\cycles[30] ),
    .C(\cycles[31] ),
    .D(_04305_),
    .X(_04309_));
 sky130_fd_sc_hd__nor2_1 _10095_ (.A(_04308_),
    .B(_04309_),
    .Y(_00028_));
 sky130_fd_sc_hd__nor2_1 _10096_ (.A(\cycles[32] ),
    .B(_04309_),
    .Y(_04310_));
 sky130_fd_sc_hd__and2_1 _10097_ (.A(\cycles[30] ),
    .B(\cycles[31] ),
    .X(_04311_));
 sky130_fd_sc_hd__and3_1 _10098_ (.A(\cycles[32] ),
    .B(_04307_),
    .C(_04311_),
    .X(_04312_));
 sky130_fd_sc_hd__nor2_1 _10099_ (.A(_04310_),
    .B(_04312_),
    .Y(_00029_));
 sky130_fd_sc_hd__and3_1 _10100_ (.A(\cycles[32] ),
    .B(\cycles[33] ),
    .C(_04309_),
    .X(_04313_));
 sky130_fd_sc_hd__o21ba_1 _10101_ (.A1(\cycles[33] ),
    .A2(_04312_),
    .B1_N(_04313_),
    .X(_00030_));
 sky130_fd_sc_hd__xor2_1 _10102_ (.A(\cycles[34] ),
    .B(_04313_),
    .X(_00031_));
 sky130_fd_sc_hd__and2_1 _10103_ (.A(\cycles[32] ),
    .B(\cycles[33] ),
    .X(_04314_));
 sky130_fd_sc_hd__and4_1 _10104_ (.A(\cycles[34] ),
    .B(_04307_),
    .C(_04311_),
    .D(_04314_),
    .X(_04315_));
 sky130_fd_sc_hd__nor2_1 _10105_ (.A(\cycles[35] ),
    .B(_04315_),
    .Y(_04316_));
 sky130_fd_sc_hd__and2_1 _10106_ (.A(\cycles[35] ),
    .B(_04315_),
    .X(_04317_));
 sky130_fd_sc_hd__nor2_1 _10107_ (.A(_04316_),
    .B(_04317_),
    .Y(_00032_));
 sky130_fd_sc_hd__nor2_1 _10108_ (.A(\cycles[36] ),
    .B(_04317_),
    .Y(_04318_));
 sky130_fd_sc_hd__and3_1 _10109_ (.A(\cycles[35] ),
    .B(\cycles[36] ),
    .C(_04315_),
    .X(_04319_));
 sky130_fd_sc_hd__nor2_1 _10110_ (.A(_04318_),
    .B(_04319_),
    .Y(_00033_));
 sky130_fd_sc_hd__and2_1 _10111_ (.A(\cycles[36] ),
    .B(\cycles[37] ),
    .X(_04320_));
 sky130_fd_sc_hd__and3_1 _10112_ (.A(\cycles[35] ),
    .B(_04315_),
    .C(_04320_),
    .X(_04321_));
 sky130_fd_sc_hd__o21ba_1 _10113_ (.A1(\cycles[37] ),
    .A2(_04319_),
    .B1_N(_04321_),
    .X(_00034_));
 sky130_fd_sc_hd__nor2_1 _10114_ (.A(\cycles[38] ),
    .B(_04321_),
    .Y(_04322_));
 sky130_fd_sc_hd__and3_1 _10115_ (.A(\cycles[34] ),
    .B(\cycles[35] ),
    .C(_04313_),
    .X(_04323_));
 sky130_fd_sc_hd__and3_1 _10116_ (.A(\cycles[38] ),
    .B(_04323_),
    .C(_04320_),
    .X(_04324_));
 sky130_fd_sc_hd__nor2_1 _10117_ (.A(_04322_),
    .B(_04324_),
    .Y(_00035_));
 sky130_fd_sc_hd__nor2_1 _10118_ (.A(\cycles[39] ),
    .B(_04324_),
    .Y(_04325_));
 sky130_fd_sc_hd__and3_1 _10119_ (.A(\cycles[38] ),
    .B(\cycles[39] ),
    .C(_04320_),
    .X(_04326_));
 sky130_fd_sc_hd__and3_1 _10120_ (.A(\cycles[35] ),
    .B(_04315_),
    .C(_04326_),
    .X(_04327_));
 sky130_fd_sc_hd__nor2_1 _10121_ (.A(_04325_),
    .B(_04327_),
    .Y(_00036_));
 sky130_fd_sc_hd__xor2_1 _10122_ (.A(\cycles[40] ),
    .B(_04327_),
    .X(_00038_));
 sky130_fd_sc_hd__a21oi_1 _10123_ (.A1(\cycles[40] ),
    .A2(_04327_),
    .B1(\cycles[41] ),
    .Y(_04328_));
 sky130_fd_sc_hd__and2_1 _10124_ (.A(\cycles[40] ),
    .B(\cycles[41] ),
    .X(_04329_));
 sky130_fd_sc_hd__and2_1 _10125_ (.A(_04327_),
    .B(_04329_),
    .X(_04330_));
 sky130_fd_sc_hd__nor2_1 _10126_ (.A(_04328_),
    .B(_04330_),
    .Y(_00039_));
 sky130_fd_sc_hd__xor2_1 _10127_ (.A(\cycles[42] ),
    .B(_04330_),
    .X(_00040_));
 sky130_fd_sc_hd__and4_1 _10128_ (.A(\cycles[39] ),
    .B(\cycles[42] ),
    .C(_04324_),
    .D(_04329_),
    .X(_04331_));
 sky130_fd_sc_hd__nor2_1 _10129_ (.A(\cycles[43] ),
    .B(_04331_),
    .Y(_04332_));
 sky130_fd_sc_hd__and3_1 _10130_ (.A(\cycles[42] ),
    .B(\cycles[43] ),
    .C(_04329_),
    .X(_04333_));
 sky130_fd_sc_hd__and4_1 _10131_ (.A(\cycles[35] ),
    .B(_04315_),
    .C(_04326_),
    .D(_04333_),
    .X(_04334_));
 sky130_fd_sc_hd__nor2_1 _10132_ (.A(_04332_),
    .B(_04334_),
    .Y(_00041_));
 sky130_fd_sc_hd__xor2_1 _10133_ (.A(\cycles[44] ),
    .B(_04334_),
    .X(_00042_));
 sky130_fd_sc_hd__a21oi_1 _10134_ (.A1(\cycles[44] ),
    .A2(_04334_),
    .B1(\cycles[45] ),
    .Y(_04335_));
 sky130_fd_sc_hd__and2_1 _10135_ (.A(\cycles[44] ),
    .B(\cycles[45] ),
    .X(_04336_));
 sky130_fd_sc_hd__and2_1 _10136_ (.A(_04334_),
    .B(_04336_),
    .X(_04337_));
 sky130_fd_sc_hd__nor2_1 _10137_ (.A(_04335_),
    .B(_04337_),
    .Y(_00043_));
 sky130_fd_sc_hd__nor2_1 _10138_ (.A(\cycles[46] ),
    .B(_04337_),
    .Y(_04338_));
 sky130_fd_sc_hd__and4_1 _10139_ (.A(\cycles[43] ),
    .B(\cycles[46] ),
    .C(_04331_),
    .D(_04336_),
    .X(_04339_));
 sky130_fd_sc_hd__nor2_1 _10140_ (.A(_04338_),
    .B(_04339_),
    .Y(_00044_));
 sky130_fd_sc_hd__xor2_1 _10141_ (.A(\cycles[47] ),
    .B(_04339_),
    .X(_00045_));
 sky130_fd_sc_hd__and4_1 _10142_ (.A(\cycles[46] ),
    .B(\cycles[47] ),
    .C(_04334_),
    .D(_04336_),
    .X(_04340_));
 sky130_fd_sc_hd__xor2_1 _10143_ (.A(\cycles[48] ),
    .B(_04340_),
    .X(_00046_));
 sky130_fd_sc_hd__a21oi_1 _10144_ (.A1(\cycles[48] ),
    .A2(_04340_),
    .B1(\cycles[49] ),
    .Y(_04341_));
 sky130_fd_sc_hd__and2_1 _10145_ (.A(\cycles[48] ),
    .B(\cycles[49] ),
    .X(_04342_));
 sky130_fd_sc_hd__and3_1 _10146_ (.A(\cycles[47] ),
    .B(_04339_),
    .C(_04342_),
    .X(_04343_));
 sky130_fd_sc_hd__nor2_1 _10147_ (.A(_04341_),
    .B(_04343_),
    .Y(_00047_));
 sky130_fd_sc_hd__xor2_1 _10148_ (.A(\cycles[50] ),
    .B(_04343_),
    .X(_00049_));
 sky130_fd_sc_hd__a21oi_1 _10149_ (.A1(\cycles[50] ),
    .A2(_04343_),
    .B1(\cycles[51] ),
    .Y(_04344_));
 sky130_fd_sc_hd__and4_1 _10150_ (.A(\cycles[50] ),
    .B(\cycles[51] ),
    .C(_04340_),
    .D(_04342_),
    .X(_04345_));
 sky130_fd_sc_hd__nor2_1 _10151_ (.A(_04344_),
    .B(_04345_),
    .Y(_00050_));
 sky130_fd_sc_hd__xor2_1 _10152_ (.A(\cycles[52] ),
    .B(_04345_),
    .X(_00051_));
 sky130_fd_sc_hd__a21oi_1 _10153_ (.A1(\cycles[52] ),
    .A2(_04345_),
    .B1(\cycles[53] ),
    .Y(_04346_));
 sky130_fd_sc_hd__and3_1 _10154_ (.A(\cycles[52] ),
    .B(\cycles[53] ),
    .C(_04345_),
    .X(_04347_));
 sky130_fd_sc_hd__nor2_1 _10155_ (.A(_04346_),
    .B(_04347_),
    .Y(_00052_));
 sky130_fd_sc_hd__xor2_1 _10156_ (.A(\cycles[54] ),
    .B(_04347_),
    .X(_00053_));
 sky130_fd_sc_hd__a21oi_1 _10157_ (.A1(\cycles[54] ),
    .A2(_04347_),
    .B1(\cycles[55] ),
    .Y(_04348_));
 sky130_fd_sc_hd__and3_1 _10158_ (.A(\cycles[54] ),
    .B(\cycles[55] ),
    .C(_04347_),
    .X(_04349_));
 sky130_fd_sc_hd__nor2_1 _10159_ (.A(_04348_),
    .B(_04349_),
    .Y(_00054_));
 sky130_fd_sc_hd__xor2_1 _10160_ (.A(\cycles[56] ),
    .B(_04349_),
    .X(_00055_));
 sky130_fd_sc_hd__a21oi_1 _10161_ (.A1(\cycles[56] ),
    .A2(_04349_),
    .B1(\cycles[57] ),
    .Y(_04350_));
 sky130_fd_sc_hd__and3_1 _10162_ (.A(\cycles[56] ),
    .B(\cycles[57] ),
    .C(_04349_),
    .X(_04351_));
 sky130_fd_sc_hd__nor2_1 _10163_ (.A(_04350_),
    .B(_04351_),
    .Y(_00056_));
 sky130_fd_sc_hd__xor2_1 _10164_ (.A(\cycles[58] ),
    .B(_04351_),
    .X(_00057_));
 sky130_fd_sc_hd__a21oi_1 _10165_ (.A1(\cycles[58] ),
    .A2(_04351_),
    .B1(\cycles[59] ),
    .Y(_04352_));
 sky130_fd_sc_hd__and3_1 _10166_ (.A(\cycles[58] ),
    .B(\cycles[59] ),
    .C(_04351_),
    .X(_04353_));
 sky130_fd_sc_hd__nor2_1 _10167_ (.A(_04352_),
    .B(_04353_),
    .Y(_00058_));
 sky130_fd_sc_hd__xor2_1 _10168_ (.A(\cycles[60] ),
    .B(_04353_),
    .X(_00060_));
 sky130_fd_sc_hd__a21oi_1 _10169_ (.A1(\cycles[60] ),
    .A2(_04353_),
    .B1(\cycles[61] ),
    .Y(_04354_));
 sky130_fd_sc_hd__and3_1 _10170_ (.A(\cycles[60] ),
    .B(\cycles[61] ),
    .C(_04353_),
    .X(_04355_));
 sky130_fd_sc_hd__nor2_1 _10171_ (.A(_04354_),
    .B(_04355_),
    .Y(_00061_));
 sky130_fd_sc_hd__or2_1 _10172_ (.A(\cycles[62] ),
    .B(_04355_),
    .X(_04356_));
 sky130_fd_sc_hd__nand2_1 _10173_ (.A(\cycles[62] ),
    .B(_04355_),
    .Y(_04357_));
 sky130_fd_sc_hd__and2_1 _10174_ (.A(_04356_),
    .B(_04357_),
    .X(_04358_));
 sky130_fd_sc_hd__clkbuf_1 _10175_ (.A(_04358_),
    .X(_00062_));
 sky130_fd_sc_hd__xnor2_1 _10176_ (.A(\cycles[63] ),
    .B(_04357_),
    .Y(_00063_));
 sky130_fd_sc_hd__nand4b_1 _10177_ (.A_N(\instr[3] ),
    .B(\instr[2] ),
    .C(\instr[1] ),
    .D(\instr[0] ),
    .Y(_04359_));
 sky130_fd_sc_hd__nand3b_4 _10178_ (.A_N(\instr[6] ),
    .B(\instr[5] ),
    .C(_01530_),
    .Y(_04360_));
 sky130_fd_sc_hd__nor2_1 _10179_ (.A(_04359_),
    .B(_04360_),
    .Y(_04361_));
 sky130_fd_sc_hd__and3_2 _10180_ (.A(_01530_),
    .B(_01854_),
    .C(_04040_),
    .X(_04362_));
 sky130_fd_sc_hd__buf_4 _10181_ (.A(_04362_),
    .X(_04363_));
 sky130_fd_sc_hd__nor2_4 _10182_ (.A(_04045_),
    .B(_04360_),
    .Y(_04364_));
 sky130_fd_sc_hd__buf_4 _10183_ (.A(_04364_),
    .X(_04365_));
 sky130_fd_sc_hd__or2_4 _10184_ (.A(_04363_),
    .B(_04365_),
    .X(_04366_));
 sky130_fd_sc_hd__nand4_1 _10185_ (.A(\instr[6] ),
    .B(\instr[5] ),
    .C(_01530_),
    .D(_01854_),
    .Y(_04367_));
 sky130_fd_sc_hd__or3b_1 _10186_ (.A(_04361_),
    .B(_04366_),
    .C_N(_04367_),
    .X(_04368_));
 sky130_fd_sc_hd__nand2_1 _10187_ (.A(_01530_),
    .B(_04040_),
    .Y(_04369_));
 sky130_fd_sc_hd__nor2_1 _10188_ (.A(_04359_),
    .B(_04369_),
    .Y(_04370_));
 sky130_fd_sc_hd__or2_1 _10189_ (.A(_01532_),
    .B(_04370_),
    .X(_04371_));
 sky130_fd_sc_hd__o21ai_2 _10190_ (.A1(_04368_),
    .A2(_04371_),
    .B1(\core_state[1] ),
    .Y(_04372_));
 sky130_fd_sc_hd__inv_2 _10191_ (.A(_04372_),
    .Y(_04373_));
 sky130_fd_sc_hd__nor2_2 _10192_ (.A(_04173_),
    .B(_04367_),
    .Y(_04374_));
 sky130_fd_sc_hd__clkbuf_4 _10193_ (.A(_04374_),
    .X(_04375_));
 sky130_fd_sc_hd__clkbuf_4 _10194_ (.A(_04375_),
    .X(_04376_));
 sky130_fd_sc_hd__nand2_1 _10195_ (.A(\B_type_imm[12] ),
    .B(_01602_),
    .Y(_04377_));
 sky130_fd_sc_hd__or2_1 _10196_ (.A(_01897_),
    .B(_04377_),
    .X(_04378_));
 sky130_fd_sc_hd__or4_1 _10197_ (.A(_01567_),
    .B(_01917_),
    .C(_01900_),
    .D(_04378_),
    .X(_04379_));
 sky130_fd_sc_hd__or3b_2 _10198_ (.A(_01564_),
    .B(_04379_),
    .C_N(_02275_),
    .X(_04380_));
 sky130_fd_sc_hd__or3_2 _10199_ (.A(_01887_),
    .B(_01595_),
    .C(_01890_),
    .X(_04381_));
 sky130_fd_sc_hd__or2_1 _10200_ (.A(_01892_),
    .B(_04381_),
    .X(_04382_));
 sky130_fd_sc_hd__nor2_2 _10201_ (.A(_04380_),
    .B(_04382_),
    .Y(_04383_));
 sky130_fd_sc_hd__clkbuf_4 _10202_ (.A(_04383_),
    .X(_04384_));
 sky130_fd_sc_hd__clkbuf_4 _10203_ (.A(_04384_),
    .X(_04385_));
 sky130_fd_sc_hd__or2_1 _10204_ (.A(_02275_),
    .B(_04379_),
    .X(_04386_));
 sky130_fd_sc_hd__or4b_2 _10205_ (.A(_01595_),
    .B(_01890_),
    .C(_01892_),
    .D_N(_01887_),
    .X(_04387_));
 sky130_fd_sc_hd__nor2_2 _10206_ (.A(_04386_),
    .B(_04387_),
    .Y(_04388_));
 sky130_fd_sc_hd__clkbuf_4 _10207_ (.A(_04388_),
    .X(_04389_));
 sky130_fd_sc_hd__clkbuf_4 _10208_ (.A(_04389_),
    .X(_04390_));
 sky130_fd_sc_hd__nor2_2 _10209_ (.A(_04382_),
    .B(_04386_),
    .Y(_04391_));
 sky130_fd_sc_hd__clkbuf_4 _10210_ (.A(_04391_),
    .X(_04392_));
 sky130_fd_sc_hd__clkbuf_4 _10211_ (.A(_04392_),
    .X(_04393_));
 sky130_fd_sc_hd__nor2_2 _10212_ (.A(_04380_),
    .B(_04387_),
    .Y(_04394_));
 sky130_fd_sc_hd__clkbuf_4 _10213_ (.A(_04394_),
    .X(_04395_));
 sky130_fd_sc_hd__nand4_1 _10214_ (.A(_01567_),
    .B(_01917_),
    .C(_01892_),
    .D(_01900_),
    .Y(_04396_));
 sky130_fd_sc_hd__or4b_1 _10215_ (.A(_02275_),
    .B(_04396_),
    .C(_01564_),
    .D_N(net35),
    .X(_04397_));
 sky130_fd_sc_hd__nor3_2 _10216_ (.A(_04381_),
    .B(_04378_),
    .C(_04397_),
    .Y(_04398_));
 sky130_fd_sc_hd__a221o_1 _10217_ (.A1(\cycles[0] ),
    .A2(_04393_),
    .B1(_04395_),
    .B2(\instret[32] ),
    .C1(_04398_),
    .X(_04399_));
 sky130_fd_sc_hd__a221o_1 _10218_ (.A1(\instret[0] ),
    .A2(_04385_),
    .B1(_04390_),
    .B2(\cycles[32] ),
    .C1(_04399_),
    .X(_04400_));
 sky130_fd_sc_hd__nand2_4 _10219_ (.A(_01688_),
    .B(_01828_),
    .Y(_04401_));
 sky130_fd_sc_hd__clkbuf_4 _10220_ (.A(_04401_),
    .X(_04402_));
 sky130_fd_sc_hd__mux2_2 _10221_ (.A0(\B_type_imm[7] ),
    .A1(\rs2_content[7] ),
    .S(_04364_),
    .X(_04403_));
 sky130_fd_sc_hd__and2_1 _10222_ (.A(_01766_),
    .B(_04403_),
    .X(_04404_));
 sky130_fd_sc_hd__inv_2 _10223_ (.A(_04404_),
    .Y(_04405_));
 sky130_fd_sc_hd__mux2_1 _10224_ (.A0(\B_type_imm[5] ),
    .A1(\rs2_content[5] ),
    .S(_04365_),
    .X(_04406_));
 sky130_fd_sc_hd__nand2_2 _10225_ (.A(_01763_),
    .B(_04406_),
    .Y(_04407_));
 sky130_fd_sc_hd__and3b_2 _10226_ (.A_N(\instr[6] ),
    .B(\instr[5] ),
    .C(\instr[4] ),
    .X(_04408_));
 sky130_fd_sc_hd__a21o_1 _10227_ (.A1(_01854_),
    .A2(_04408_),
    .B1(\I_type_imm[3] ),
    .X(_04409_));
 sky130_fd_sc_hd__or3_1 _10228_ (.A(\rs2_content[3] ),
    .B(_04045_),
    .C(_04360_),
    .X(_04410_));
 sky130_fd_sc_hd__and2_1 _10229_ (.A(_04409_),
    .B(_04410_),
    .X(_04411_));
 sky130_fd_sc_hd__nand2_1 _10230_ (.A(_01771_),
    .B(_04411_),
    .Y(_04412_));
 sky130_fd_sc_hd__a21o_1 _10231_ (.A1(_01854_),
    .A2(_04408_),
    .B1(\I_type_imm[1] ),
    .X(_04413_));
 sky130_fd_sc_hd__or3_1 _10232_ (.A(\rs2_content[1] ),
    .B(_04045_),
    .C(_04360_),
    .X(_04414_));
 sky130_fd_sc_hd__and3_1 _10233_ (.A(\leorv32_alu.input1[1] ),
    .B(_04413_),
    .C(_04414_),
    .X(_04415_));
 sky130_fd_sc_hd__a21oi_1 _10234_ (.A1(_04413_),
    .A2(_04414_),
    .B1(_01778_),
    .Y(_04416_));
 sky130_fd_sc_hd__nor2_1 _10235_ (.A(_04415_),
    .B(_04416_),
    .Y(_04417_));
 sky130_fd_sc_hd__mux2_1 _10236_ (.A0(\I_type_imm[0] ),
    .A1(\rs2_content[0] ),
    .S(_04364_),
    .X(_04418_));
 sky130_fd_sc_hd__nor2_1 _10237_ (.A(_01807_),
    .B(_04418_),
    .Y(_04419_));
 sky130_fd_sc_hd__and2_1 _10238_ (.A(_01807_),
    .B(_04418_),
    .X(_04420_));
 sky130_fd_sc_hd__nor2_1 _10239_ (.A(_04419_),
    .B(_04420_),
    .Y(_04421_));
 sky130_fd_sc_hd__and3_1 _10240_ (.A(\leorv32_alu.input1[3] ),
    .B(_04409_),
    .C(_04410_),
    .X(_04422_));
 sky130_fd_sc_hd__a21oi_1 _10241_ (.A1(_04409_),
    .A2(_04410_),
    .B1(_01898_),
    .Y(_04423_));
 sky130_fd_sc_hd__nor2_2 _10242_ (.A(_04422_),
    .B(_04423_),
    .Y(_04424_));
 sky130_fd_sc_hd__inv_2 _10243_ (.A(\I_type_imm[2] ),
    .Y(_04425_));
 sky130_fd_sc_hd__inv_2 _10244_ (.A(\rs2_content[2] ),
    .Y(_04426_));
 sky130_fd_sc_hd__mux2_2 _10245_ (.A0(_04425_),
    .A1(_04426_),
    .S(_04364_),
    .X(_04427_));
 sky130_fd_sc_hd__xnor2_2 _10246_ (.A(\leorv32_alu.input1[2] ),
    .B(_04427_),
    .Y(_04428_));
 sky130_fd_sc_hd__or4_1 _10247_ (.A(_04417_),
    .B(_04421_),
    .C(_04424_),
    .D(_04428_),
    .X(_04429_));
 sky130_fd_sc_hd__a2bb2o_1 _10248_ (.A1_N(_04415_),
    .A2_N(_04416_),
    .B1(_04418_),
    .B2(_01776_),
    .X(_04430_));
 sky130_fd_sc_hd__a21o_1 _10249_ (.A1(_04413_),
    .A2(_04414_),
    .B1(_01775_),
    .X(_04431_));
 sky130_fd_sc_hd__a21oi_1 _10250_ (.A1(_04430_),
    .A2(_04431_),
    .B1(_04428_),
    .Y(_04432_));
 sky130_fd_sc_hd__a21oi_1 _10251_ (.A1(_01901_),
    .A2(_04427_),
    .B1(_04432_),
    .Y(_04433_));
 sky130_fd_sc_hd__o21ai_1 _10252_ (.A1(_01771_),
    .A2(_04411_),
    .B1(_04433_),
    .Y(_04434_));
 sky130_fd_sc_hd__mux2_1 _10253_ (.A0(\I_type_imm[4] ),
    .A1(\rs2_content[4] ),
    .S(_04365_),
    .X(_04435_));
 sky130_fd_sc_hd__and2_2 _10254_ (.A(\leorv32_alu.input1[4] ),
    .B(_04435_),
    .X(_04436_));
 sky130_fd_sc_hd__nor2_1 _10255_ (.A(_01764_),
    .B(_04435_),
    .Y(_04437_));
 sky130_fd_sc_hd__nor2_2 _10256_ (.A(_04436_),
    .B(_04437_),
    .Y(_04438_));
 sky130_fd_sc_hd__a31o_1 _10257_ (.A1(_04412_),
    .A2(_04429_),
    .A3(_04434_),
    .B1(_04438_),
    .X(_04439_));
 sky130_fd_sc_hd__nand2_1 _10258_ (.A(_01765_),
    .B(_04435_),
    .Y(_04440_));
 sky130_fd_sc_hd__or2_1 _10259_ (.A(_01763_),
    .B(_04406_),
    .X(_04441_));
 sky130_fd_sc_hd__inv_2 _10260_ (.A(_04441_),
    .Y(_04442_));
 sky130_fd_sc_hd__xnor2_2 _10261_ (.A(_01766_),
    .B(_04403_),
    .Y(_04443_));
 sky130_fd_sc_hd__mux2_2 _10262_ (.A0(\B_type_imm[6] ),
    .A1(\rs2_content[6] ),
    .S(_04364_),
    .X(_04444_));
 sky130_fd_sc_hd__xnor2_2 _10263_ (.A(_01767_),
    .B(_04444_),
    .Y(_04445_));
 sky130_fd_sc_hd__or2_1 _10264_ (.A(_04443_),
    .B(_04445_),
    .X(_04446_));
 sky130_fd_sc_hd__a311o_1 _10265_ (.A1(_04407_),
    .A2(_04439_),
    .A3(_04440_),
    .B1(_04442_),
    .C1(_04446_),
    .X(_04447_));
 sky130_fd_sc_hd__or2_1 _10266_ (.A(_01766_),
    .B(_04403_),
    .X(_04448_));
 sky130_fd_sc_hd__nand3_1 _10267_ (.A(_01767_),
    .B(_04448_),
    .C(_04444_),
    .Y(_04449_));
 sky130_fd_sc_hd__nand2_1 _10268_ (.A(_01854_),
    .B(_04408_),
    .Y(_04450_));
 sky130_fd_sc_hd__a21o_1 _10269_ (.A1(_01854_),
    .A2(_04408_),
    .B1(\B_type_imm[12] ),
    .X(_04451_));
 sky130_fd_sc_hd__o21a_2 _10270_ (.A1(\rs2_content[15] ),
    .A2(_04450_),
    .B1(_04451_),
    .X(_04452_));
 sky130_fd_sc_hd__xor2_2 _10271_ (.A(\leorv32_alu.input1[15] ),
    .B(_04452_),
    .X(_04453_));
 sky130_fd_sc_hd__buf_2 _10272_ (.A(_04451_),
    .X(_04454_));
 sky130_fd_sc_hd__or3_1 _10273_ (.A(\rs2_content[14] ),
    .B(_04045_),
    .C(_04360_),
    .X(_04455_));
 sky130_fd_sc_hd__and3_1 _10274_ (.A(\leorv32_alu.input1[14] ),
    .B(_04454_),
    .C(_04455_),
    .X(_04456_));
 sky130_fd_sc_hd__a21oi_1 _10275_ (.A1(_04454_),
    .A2(_04455_),
    .B1(_01871_),
    .Y(_04457_));
 sky130_fd_sc_hd__nor2_1 _10276_ (.A(_04456_),
    .B(_04457_),
    .Y(_04458_));
 sky130_fd_sc_hd__or2_1 _10277_ (.A(_04453_),
    .B(_04458_),
    .X(_04459_));
 sky130_fd_sc_hd__clkbuf_4 _10278_ (.A(_04450_),
    .X(_04460_));
 sky130_fd_sc_hd__o21a_1 _10279_ (.A1(\rs2_content[13] ),
    .A2(_04460_),
    .B1(_04454_),
    .X(_04461_));
 sky130_fd_sc_hd__or2b_1 _10280_ (.A(_04461_),
    .B_N(_01872_),
    .X(_04462_));
 sky130_fd_sc_hd__nand2b_2 _10281_ (.A_N(\leorv32_alu.input1[13] ),
    .B(_04461_),
    .Y(_04463_));
 sky130_fd_sc_hd__nand2_1 _10282_ (.A(_04462_),
    .B(_04463_),
    .Y(_04464_));
 sky130_fd_sc_hd__o211a_1 _10283_ (.A1(\rs2_content[12] ),
    .A2(_04460_),
    .B1(_04454_),
    .C1(\leorv32_alu.input1[12] ),
    .X(_04465_));
 sky130_fd_sc_hd__o21ai_1 _10284_ (.A1(\rs2_content[12] ),
    .A2(_04460_),
    .B1(_04454_),
    .Y(_04466_));
 sky130_fd_sc_hd__and2b_1 _10285_ (.A_N(\leorv32_alu.input1[12] ),
    .B(_04466_),
    .X(_04467_));
 sky130_fd_sc_hd__or2_1 _10286_ (.A(_04465_),
    .B(_04467_),
    .X(_04468_));
 sky130_fd_sc_hd__or3b_1 _10287_ (.A(_04459_),
    .B(_04464_),
    .C_N(_04468_),
    .X(_04469_));
 sky130_fd_sc_hd__mux2_1 _10288_ (.A0(_01879_),
    .A1(_01750_),
    .S(_04364_),
    .X(_04470_));
 sky130_fd_sc_hd__nor2_2 _10289_ (.A(_01880_),
    .B(_04470_),
    .Y(_04471_));
 sky130_fd_sc_hd__mux2_1 _10290_ (.A0(\barrel_shifter_right.arith ),
    .A1(\rs2_content[10] ),
    .S(_04365_),
    .X(_04472_));
 sky130_fd_sc_hd__nor2_1 _10291_ (.A(_01877_),
    .B(_04472_),
    .Y(_04473_));
 sky130_fd_sc_hd__nor2_2 _10292_ (.A(_04471_),
    .B(_04473_),
    .Y(_04474_));
 sky130_fd_sc_hd__o21ai_1 _10293_ (.A1(\rs2_content[11] ),
    .A2(_04460_),
    .B1(_04454_),
    .Y(_04475_));
 sky130_fd_sc_hd__and2_1 _10294_ (.A(\leorv32_alu.input1[11] ),
    .B(_04475_),
    .X(_04476_));
 sky130_fd_sc_hd__or2_2 _10295_ (.A(\leorv32_alu.input1[11] ),
    .B(_04475_),
    .X(_04477_));
 sky130_fd_sc_hd__nand2b_2 _10296_ (.A_N(_04476_),
    .B(_04477_),
    .Y(_04478_));
 sky130_fd_sc_hd__or2_1 _10297_ (.A(_04474_),
    .B(_04478_),
    .X(_04479_));
 sky130_fd_sc_hd__mux2_2 _10298_ (.A0(\B_type_imm[8] ),
    .A1(\rs2_content[8] ),
    .S(_04365_),
    .X(_04480_));
 sky130_fd_sc_hd__and2_1 _10299_ (.A(\leorv32_alu.input1[8] ),
    .B(_04480_),
    .X(_04481_));
 sky130_fd_sc_hd__nor2_1 _10300_ (.A(\leorv32_alu.input1[8] ),
    .B(_04480_),
    .Y(_04482_));
 sky130_fd_sc_hd__nor2_2 _10301_ (.A(_04481_),
    .B(_04482_),
    .Y(_04483_));
 sky130_fd_sc_hd__inv_2 _10302_ (.A(_01752_),
    .Y(_04484_));
 sky130_fd_sc_hd__mux2_2 _10303_ (.A0(\B_type_imm[9] ),
    .A1(\rs2_content[9] ),
    .S(_04365_),
    .X(_04485_));
 sky130_fd_sc_hd__and2_1 _10304_ (.A(_04484_),
    .B(_04485_),
    .X(_04486_));
 sky130_fd_sc_hd__nor2_1 _10305_ (.A(_04484_),
    .B(_04485_),
    .Y(_04487_));
 sky130_fd_sc_hd__or2_2 _10306_ (.A(_04486_),
    .B(_04487_),
    .X(_04488_));
 sky130_fd_sc_hd__or4_2 _10307_ (.A(_04469_),
    .B(_04479_),
    .C(_04483_),
    .D(_04488_),
    .X(_04489_));
 sky130_fd_sc_hd__a31o_1 _10308_ (.A1(_04405_),
    .A2(_04447_),
    .A3(_04449_),
    .B1(_04489_),
    .X(_04490_));
 sky130_fd_sc_hd__a21oi_1 _10309_ (.A1(_01754_),
    .A2(_04480_),
    .B1(_04486_),
    .Y(_04491_));
 sky130_fd_sc_hd__or3_1 _10310_ (.A(_01877_),
    .B(_04470_),
    .C(_04476_),
    .X(_04492_));
 sky130_fd_sc_hd__o311a_1 _10311_ (.A1(_04479_),
    .A2(_04487_),
    .A3(_04491_),
    .B1(_04492_),
    .C1(_04477_),
    .X(_04493_));
 sky130_fd_sc_hd__and2b_1 _10312_ (.A_N(_04461_),
    .B(_01872_),
    .X(_04494_));
 sky130_fd_sc_hd__o31a_1 _10313_ (.A1(_01747_),
    .A2(_04494_),
    .A3(_04466_),
    .B1(_04463_),
    .X(_04495_));
 sky130_fd_sc_hd__and2b_1 _10314_ (.A_N(_04452_),
    .B(_01870_),
    .X(_04496_));
 sky130_fd_sc_hd__buf_2 _10315_ (.A(_04454_),
    .X(_04497_));
 sky130_fd_sc_hd__clkbuf_4 _10316_ (.A(_04497_),
    .X(_04498_));
 sky130_fd_sc_hd__nand2_1 _10317_ (.A(_04498_),
    .B(_04455_),
    .Y(_04499_));
 sky130_fd_sc_hd__or2b_1 _10318_ (.A(_01870_),
    .B_N(_04452_),
    .X(_04500_));
 sky130_fd_sc_hd__o31a_1 _10319_ (.A1(_01871_),
    .A2(_04496_),
    .A3(_04499_),
    .B1(_04500_),
    .X(_04501_));
 sky130_fd_sc_hd__o221a_1 _10320_ (.A1(_04469_),
    .A2(_04493_),
    .B1(_04495_),
    .B2(_04459_),
    .C1(_04501_),
    .X(_04502_));
 sky130_fd_sc_hd__clkbuf_4 _10321_ (.A(_04460_),
    .X(_04503_));
 sky130_fd_sc_hd__o21a_1 _10322_ (.A1(\rs2_content[18] ),
    .A2(_04503_),
    .B1(_04497_),
    .X(_04504_));
 sky130_fd_sc_hd__and2_1 _10323_ (.A(_01867_),
    .B(_04504_),
    .X(_04505_));
 sky130_fd_sc_hd__nor2_1 _10324_ (.A(_01867_),
    .B(_04504_),
    .Y(_04506_));
 sky130_fd_sc_hd__or2_1 _10325_ (.A(_04505_),
    .B(_04506_),
    .X(_04507_));
 sky130_fd_sc_hd__inv_2 _10326_ (.A(_01717_),
    .Y(_04508_));
 sky130_fd_sc_hd__o21a_1 _10327_ (.A1(\rs2_content[19] ),
    .A2(_04460_),
    .B1(_04497_),
    .X(_04509_));
 sky130_fd_sc_hd__or2_1 _10328_ (.A(_04508_),
    .B(_04509_),
    .X(_04510_));
 sky130_fd_sc_hd__inv_2 _10329_ (.A(_04510_),
    .Y(_04511_));
 sky130_fd_sc_hd__and2_1 _10330_ (.A(_04508_),
    .B(_04509_),
    .X(_04512_));
 sky130_fd_sc_hd__nor2_1 _10331_ (.A(_04511_),
    .B(_04512_),
    .Y(_04513_));
 sky130_fd_sc_hd__nand2_1 _10332_ (.A(_04507_),
    .B(_04513_),
    .Y(_04514_));
 sky130_fd_sc_hd__inv_2 _10333_ (.A(_01723_),
    .Y(_04515_));
 sky130_fd_sc_hd__o21a_1 _10334_ (.A1(\rs2_content[17] ),
    .A2(_04503_),
    .B1(_04497_),
    .X(_04516_));
 sky130_fd_sc_hd__or2_1 _10335_ (.A(_04515_),
    .B(_04516_),
    .X(_04517_));
 sky130_fd_sc_hd__nand2_1 _10336_ (.A(_04515_),
    .B(_04516_),
    .Y(_04518_));
 sky130_fd_sc_hd__nand2_2 _10337_ (.A(_04517_),
    .B(_04518_),
    .Y(_04519_));
 sky130_fd_sc_hd__buf_4 _10338_ (.A(_04503_),
    .X(_04520_));
 sky130_fd_sc_hd__o21ai_2 _10339_ (.A1(\rs2_content[16] ),
    .A2(_04520_),
    .B1(_04498_),
    .Y(_04521_));
 sky130_fd_sc_hd__nor2_2 _10340_ (.A(_01799_),
    .B(_04521_),
    .Y(_04522_));
 sky130_fd_sc_hd__o21a_1 _10341_ (.A1(\rs2_content[16] ),
    .A2(_04503_),
    .B1(_04498_),
    .X(_04523_));
 sky130_fd_sc_hd__nor2_1 _10342_ (.A(_01868_),
    .B(_04523_),
    .Y(_04524_));
 sky130_fd_sc_hd__nor2_2 _10343_ (.A(_04522_),
    .B(_04524_),
    .Y(_04525_));
 sky130_fd_sc_hd__o21ai_1 _10344_ (.A1(\rs2_content[22] ),
    .A2(_04503_),
    .B1(_04497_),
    .Y(_04526_));
 sky130_fd_sc_hd__nor2_2 _10345_ (.A(_01712_),
    .B(_04526_),
    .Y(_04527_));
 sky130_fd_sc_hd__o21a_1 _10346_ (.A1(\rs2_content[22] ),
    .A2(_04503_),
    .B1(_04497_),
    .X(_04528_));
 sky130_fd_sc_hd__nor2_1 _10347_ (.A(\leorv32_alu.input1[22] ),
    .B(_04528_),
    .Y(_04529_));
 sky130_fd_sc_hd__nor2_1 _10348_ (.A(_04527_),
    .B(_04529_),
    .Y(_04530_));
 sky130_fd_sc_hd__o21a_1 _10349_ (.A1(\rs2_content[23] ),
    .A2(_04460_),
    .B1(_04454_),
    .X(_04531_));
 sky130_fd_sc_hd__or2_1 _10350_ (.A(_01711_),
    .B(_04531_),
    .X(_04532_));
 sky130_fd_sc_hd__nand2_1 _10351_ (.A(_01711_),
    .B(_04531_),
    .Y(_04533_));
 sky130_fd_sc_hd__nand2_2 _10352_ (.A(_04532_),
    .B(_04533_),
    .Y(_04534_));
 sky130_fd_sc_hd__or2_1 _10353_ (.A(_04530_),
    .B(_04534_),
    .X(_04535_));
 sky130_fd_sc_hd__o21a_1 _10354_ (.A1(\rs2_content[21] ),
    .A2(_04460_),
    .B1(_04454_),
    .X(_04536_));
 sky130_fd_sc_hd__and2_1 _10355_ (.A(\leorv32_alu.input1[21] ),
    .B(_04536_),
    .X(_04537_));
 sky130_fd_sc_hd__inv_2 _10356_ (.A(_04537_),
    .Y(_04538_));
 sky130_fd_sc_hd__or2_1 _10357_ (.A(\leorv32_alu.input1[21] ),
    .B(_04536_),
    .X(_04539_));
 sky130_fd_sc_hd__and2_2 _10358_ (.A(_04538_),
    .B(_04539_),
    .X(_04540_));
 sky130_fd_sc_hd__o21ai_2 _10359_ (.A1(\rs2_content[20] ),
    .A2(_04460_),
    .B1(_04454_),
    .Y(_04541_));
 sky130_fd_sc_hd__and2_1 _10360_ (.A(_01715_),
    .B(_04541_),
    .X(_04542_));
 sky130_fd_sc_hd__nor2_2 _10361_ (.A(_01715_),
    .B(_04541_),
    .Y(_04543_));
 sky130_fd_sc_hd__or2_1 _10362_ (.A(_04542_),
    .B(_04543_),
    .X(_04544_));
 sky130_fd_sc_hd__inv_2 _10363_ (.A(_04544_),
    .Y(_04545_));
 sky130_fd_sc_hd__or3_1 _10364_ (.A(_04535_),
    .B(_04540_),
    .C(_04545_),
    .X(_04546_));
 sky130_fd_sc_hd__or4_2 _10365_ (.A(_04514_),
    .B(_04519_),
    .C(_04525_),
    .D(_04546_),
    .X(_04547_));
 sky130_fd_sc_hd__a21o_1 _10366_ (.A1(_04490_),
    .A2(_04502_),
    .B1(_04547_),
    .X(_04548_));
 sky130_fd_sc_hd__o21a_1 _10367_ (.A1(_01868_),
    .A2(_04521_),
    .B1(_04518_),
    .X(_04549_));
 sky130_fd_sc_hd__nor2_1 _10368_ (.A(_04514_),
    .B(_04549_),
    .Y(_04550_));
 sky130_fd_sc_hd__inv_2 _10369_ (.A(_01867_),
    .Y(_04551_));
 sky130_fd_sc_hd__a31o_1 _10370_ (.A1(_04551_),
    .A2(_04504_),
    .A3(_04510_),
    .B1(_04512_),
    .X(_04552_));
 sky130_fd_sc_hd__a21oi_1 _10371_ (.A1(_04517_),
    .A2(_04550_),
    .B1(_04552_),
    .Y(_04553_));
 sky130_fd_sc_hd__nor2_1 _10372_ (.A(_01714_),
    .B(_04536_),
    .Y(_04554_));
 sky130_fd_sc_hd__nand2_1 _10373_ (.A(_01714_),
    .B(_04536_),
    .Y(_04555_));
 sky130_fd_sc_hd__o31a_1 _10374_ (.A1(\leorv32_alu.input1[20] ),
    .A2(_04554_),
    .A3(_04541_),
    .B1(_04555_),
    .X(_04556_));
 sky130_fd_sc_hd__inv_2 _10375_ (.A(_04533_),
    .Y(_04557_));
 sky130_fd_sc_hd__a31oi_1 _10376_ (.A1(_01712_),
    .A2(_04528_),
    .A3(_04532_),
    .B1(_04557_),
    .Y(_04558_));
 sky130_fd_sc_hd__o221a_1 _10377_ (.A1(_04546_),
    .A2(_04553_),
    .B1(_04556_),
    .B2(_04535_),
    .C1(_04558_),
    .X(_04559_));
 sky130_fd_sc_hd__o21a_1 _10378_ (.A1(\rs2_content[25] ),
    .A2(_04503_),
    .B1(_04497_),
    .X(_04560_));
 sky130_fd_sc_hd__and2_1 _10379_ (.A(\leorv32_alu.input1[25] ),
    .B(_04560_),
    .X(_04561_));
 sky130_fd_sc_hd__or2_1 _10380_ (.A(\leorv32_alu.input1[25] ),
    .B(_04560_),
    .X(_04562_));
 sky130_fd_sc_hd__nor2b_2 _10381_ (.A(_04561_),
    .B_N(_04562_),
    .Y(_04563_));
 sky130_fd_sc_hd__o21a_1 _10382_ (.A1(\rs2_content[24] ),
    .A2(_04520_),
    .B1(_04498_),
    .X(_04564_));
 sky130_fd_sc_hd__nor2_1 _10383_ (.A(\leorv32_alu.input1[24] ),
    .B(_04564_),
    .Y(_04565_));
 sky130_fd_sc_hd__and2_1 _10384_ (.A(\leorv32_alu.input1[24] ),
    .B(_04564_),
    .X(_04566_));
 sky130_fd_sc_hd__nor2_2 _10385_ (.A(_04565_),
    .B(_04566_),
    .Y(_04567_));
 sky130_fd_sc_hd__o21ai_2 _10386_ (.A1(\rs2_content[26] ),
    .A2(_04503_),
    .B1(_04497_),
    .Y(_04568_));
 sky130_fd_sc_hd__nor2_1 _10387_ (.A(_01705_),
    .B(_04568_),
    .Y(_04569_));
 sky130_fd_sc_hd__and2_1 _10388_ (.A(_01705_),
    .B(_04568_),
    .X(_04570_));
 sky130_fd_sc_hd__or2_2 _10389_ (.A(_04569_),
    .B(_04570_),
    .X(_04571_));
 sky130_fd_sc_hd__o21ai_2 _10390_ (.A1(\rs2_content[27] ),
    .A2(_04460_),
    .B1(_04497_),
    .Y(_04572_));
 sky130_fd_sc_hd__or2_1 _10391_ (.A(\leorv32_alu.input1[27] ),
    .B(_04572_),
    .X(_04573_));
 sky130_fd_sc_hd__nand2_1 _10392_ (.A(\leorv32_alu.input1[27] ),
    .B(_04572_),
    .Y(_04574_));
 sky130_fd_sc_hd__and2_1 _10393_ (.A(_04573_),
    .B(_04574_),
    .X(_04575_));
 sky130_fd_sc_hd__clkbuf_2 _10394_ (.A(_04575_),
    .X(_04576_));
 sky130_fd_sc_hd__and2_1 _10395_ (.A(_04571_),
    .B(_04576_),
    .X(_04577_));
 sky130_fd_sc_hd__nor3b_1 _10396_ (.A(_04563_),
    .B(_04567_),
    .C_N(_04577_),
    .Y(_04578_));
 sky130_fd_sc_hd__inv_2 _10397_ (.A(_04578_),
    .Y(_04579_));
 sky130_fd_sc_hd__o21ai_1 _10398_ (.A1(\rs2_content[29] ),
    .A2(_04520_),
    .B1(_04498_),
    .Y(_04580_));
 sky130_fd_sc_hd__or2_1 _10399_ (.A(\leorv32_alu.input1[29] ),
    .B(_04580_),
    .X(_04581_));
 sky130_fd_sc_hd__nand2_1 _10400_ (.A(\leorv32_alu.input1[29] ),
    .B(_04580_),
    .Y(_04582_));
 sky130_fd_sc_hd__nand2_2 _10401_ (.A(_04581_),
    .B(_04582_),
    .Y(_04583_));
 sky130_fd_sc_hd__o21a_1 _10402_ (.A1(\rs2_content[31] ),
    .A2(_04503_),
    .B1(_04498_),
    .X(_04584_));
 sky130_fd_sc_hd__xnor2_1 _10403_ (.A(\leorv32_alu.input1[31] ),
    .B(_04584_),
    .Y(_04585_));
 sky130_fd_sc_hd__inv_2 _10404_ (.A(_04585_),
    .Y(_04586_));
 sky130_fd_sc_hd__o21a_1 _10405_ (.A1(\rs2_content[28] ),
    .A2(_04520_),
    .B1(_04498_),
    .X(_04587_));
 sky130_fd_sc_hd__or2b_1 _10406_ (.A(_01736_),
    .B_N(_04587_),
    .X(_04588_));
 sky130_fd_sc_hd__nand2b_1 _10407_ (.A_N(_04587_),
    .B(_01736_),
    .Y(_04589_));
 sky130_fd_sc_hd__nand2_1 _10408_ (.A(_04588_),
    .B(_04589_),
    .Y(_04590_));
 sky130_fd_sc_hd__o21a_1 _10409_ (.A1(\rs2_content[30] ),
    .A2(_04520_),
    .B1(_04498_),
    .X(_04591_));
 sky130_fd_sc_hd__nor2_1 _10410_ (.A(\leorv32_alu.input1[30] ),
    .B(_04591_),
    .Y(_04592_));
 sky130_fd_sc_hd__o21ai_2 _10411_ (.A1(\rs2_content[30] ),
    .A2(_04520_),
    .B1(_04498_),
    .Y(_04593_));
 sky130_fd_sc_hd__nor2_1 _10412_ (.A(_01694_),
    .B(_04593_),
    .Y(_04594_));
 sky130_fd_sc_hd__nor2_1 _10413_ (.A(_04592_),
    .B(_04594_),
    .Y(_04595_));
 sky130_fd_sc_hd__or4_1 _10414_ (.A(_04583_),
    .B(_04586_),
    .C(_04590_),
    .D(_04595_),
    .X(_04596_));
 sky130_fd_sc_hd__or2_1 _10415_ (.A(_04579_),
    .B(_04596_),
    .X(_04597_));
 sky130_fd_sc_hd__a21o_1 _10416_ (.A1(_04548_),
    .A2(_04559_),
    .B1(_04597_),
    .X(_04598_));
 sky130_fd_sc_hd__nand2_1 _10417_ (.A(_01702_),
    .B(_04560_),
    .Y(_04599_));
 sky130_fd_sc_hd__nand2_1 _10418_ (.A(_01703_),
    .B(_04564_),
    .Y(_04600_));
 sky130_fd_sc_hd__nor2_1 _10419_ (.A(_01702_),
    .B(_04560_),
    .Y(_04601_));
 sky130_fd_sc_hd__a221o_1 _10420_ (.A1(\leorv32_alu.input1[26] ),
    .A2(_04568_),
    .B1(_04599_),
    .B2(_04600_),
    .C1(_04601_),
    .X(_04602_));
 sky130_fd_sc_hd__o211ai_1 _10421_ (.A1(\leorv32_alu.input1[26] ),
    .A2(_04568_),
    .B1(_04573_),
    .C1(_04602_),
    .Y(_04603_));
 sky130_fd_sc_hd__nand2_1 _10422_ (.A(_04581_),
    .B(_04588_),
    .Y(_04604_));
 sky130_fd_sc_hd__a31oi_1 _10423_ (.A1(_04574_),
    .A2(_04589_),
    .A3(_04603_),
    .B1(_04604_),
    .Y(_04605_));
 sky130_fd_sc_hd__o21ai_1 _10424_ (.A1(_01694_),
    .A2(_04591_),
    .B1(_04582_),
    .Y(_04606_));
 sky130_fd_sc_hd__o22a_1 _10425_ (.A1(\leorv32_alu.input1[30] ),
    .A2(_04593_),
    .B1(_04605_),
    .B2(_04606_),
    .X(_04607_));
 sky130_fd_sc_hd__or2b_1 _10426_ (.A(\leorv32_alu.input1[31] ),
    .B_N(_04584_),
    .X(_04608_));
 sky130_fd_sc_hd__o21a_1 _10427_ (.A1(_04586_),
    .A2(_04607_),
    .B1(_04608_),
    .X(_04609_));
 sky130_fd_sc_hd__nor2_1 _10428_ (.A(_01826_),
    .B(_04585_),
    .Y(_04610_));
 sky130_fd_sc_hd__a21boi_1 _10429_ (.A1(_04598_),
    .A2(_04609_),
    .B1_N(_04610_),
    .Y(_04611_));
 sky130_fd_sc_hd__nand2_2 _10430_ (.A(_04441_),
    .B(_04407_),
    .Y(_04612_));
 sky130_fd_sc_hd__or4_1 _10431_ (.A(_04446_),
    .B(_04438_),
    .C(_04612_),
    .D(_04429_),
    .X(_04613_));
 sky130_fd_sc_hd__nor4_1 _10432_ (.A(_04597_),
    .B(_04547_),
    .C(_04489_),
    .D(_04613_),
    .Y(_04614_));
 sky130_fd_sc_hd__o211a_1 _10433_ (.A1(_01826_),
    .A2(_04585_),
    .B1(_04598_),
    .C1(_04609_),
    .X(_04615_));
 sky130_fd_sc_hd__or4_1 _10434_ (.A(_01979_),
    .B(_04611_),
    .C(_04614_),
    .D(_04615_),
    .X(_04616_));
 sky130_fd_sc_hd__nor4_4 _10435_ (.A(_01535_),
    .B(_01567_),
    .C(_01917_),
    .D(_04381_),
    .Y(_04617_));
 sky130_fd_sc_hd__nor2_1 _10436_ (.A(_01688_),
    .B(_04617_),
    .Y(_04618_));
 sky130_fd_sc_hd__or2_1 _10437_ (.A(_01969_),
    .B(_04618_),
    .X(_04619_));
 sky130_fd_sc_hd__mux2_2 _10438_ (.A0(\rs2_content[1] ),
    .A1(\I_type_imm[1] ),
    .S(_04363_),
    .X(_04620_));
 sky130_fd_sc_hd__buf_2 _10439_ (.A(_04620_),
    .X(_04621_));
 sky130_fd_sc_hd__buf_2 _10440_ (.A(_04621_),
    .X(_04622_));
 sky130_fd_sc_hd__mux2_1 _10441_ (.A0(\leorv32_alu.input1[30] ),
    .A1(_01778_),
    .S(_01686_),
    .X(_04623_));
 sky130_fd_sc_hd__clkbuf_4 _10442_ (.A(\J_type_imm[14] ),
    .X(_04624_));
 sky130_fd_sc_hd__mux2_1 _10443_ (.A0(_01871_),
    .A1(_01723_),
    .S(_04624_),
    .X(_04625_));
 sky130_fd_sc_hd__mux2_4 _10444_ (.A0(\rs2_content[4] ),
    .A1(\I_type_imm[4] ),
    .S(_04362_),
    .X(_04626_));
 sky130_fd_sc_hd__buf_2 _10445_ (.A(_04626_),
    .X(_04627_));
 sky130_fd_sc_hd__clkbuf_4 _10446_ (.A(_04627_),
    .X(_04628_));
 sky130_fd_sc_hd__mux2_1 _10447_ (.A0(_04623_),
    .A1(_04625_),
    .S(_04628_),
    .X(_04629_));
 sky130_fd_sc_hd__mux2_1 _10448_ (.A0(\leorv32_alu.input1[22] ),
    .A1(_01752_),
    .S(_01686_),
    .X(_04630_));
 sky130_fd_sc_hd__mux2_1 _10449_ (.A0(\leorv32_alu.input1[6] ),
    .A1(\leorv32_alu.input1[25] ),
    .S(_04624_),
    .X(_04631_));
 sky130_fd_sc_hd__mux2_1 _10450_ (.A0(_04630_),
    .A1(_04631_),
    .S(_04628_),
    .X(_04632_));
 sky130_fd_sc_hd__mux2_4 _10451_ (.A0(_01770_),
    .A1(_01897_),
    .S(_04362_),
    .X(_04633_));
 sky130_fd_sc_hd__buf_2 _10452_ (.A(_04633_),
    .X(_04634_));
 sky130_fd_sc_hd__buf_2 _10453_ (.A(_04634_),
    .X(_04635_));
 sky130_fd_sc_hd__mux2_1 _10454_ (.A0(_04629_),
    .A1(_04632_),
    .S(_04635_),
    .X(_04636_));
 sky130_fd_sc_hd__mux2_1 _10455_ (.A0(_01867_),
    .A1(_01872_),
    .S(_01685_),
    .X(_04637_));
 sky130_fd_sc_hd__mux2_1 _10456_ (.A0(_01901_),
    .A1(\leorv32_alu.input1[29] ),
    .S(_01685_),
    .X(_04638_));
 sky130_fd_sc_hd__mux2_1 _10457_ (.A0(_04637_),
    .A1(_04638_),
    .S(_04626_),
    .X(_04639_));
 sky130_fd_sc_hd__mux2_1 _10458_ (.A0(\leorv32_alu.input1[26] ),
    .A1(\leorv32_alu.input1[5] ),
    .S(_01686_),
    .X(_04640_));
 sky130_fd_sc_hd__mux2_1 _10459_ (.A0(_01877_),
    .A1(\leorv32_alu.input1[21] ),
    .S(_04624_),
    .X(_04641_));
 sky130_fd_sc_hd__mux2_1 _10460_ (.A0(_04640_),
    .A1(_04641_),
    .S(_04628_),
    .X(_04642_));
 sky130_fd_sc_hd__inv_2 _10461_ (.A(_01770_),
    .Y(_04643_));
 sky130_fd_sc_hd__inv_2 _10462_ (.A(_01897_),
    .Y(_04644_));
 sky130_fd_sc_hd__mux2_4 _10463_ (.A0(_04643_),
    .A1(_04644_),
    .S(_04363_),
    .X(_04645_));
 sky130_fd_sc_hd__buf_2 _10464_ (.A(_04645_),
    .X(_04646_));
 sky130_fd_sc_hd__mux2_1 _10465_ (.A0(_04639_),
    .A1(_04642_),
    .S(_04646_),
    .X(_04647_));
 sky130_fd_sc_hd__mux2_4 _10466_ (.A0(_01772_),
    .A1(_01900_),
    .S(_04363_),
    .X(_04648_));
 sky130_fd_sc_hd__buf_2 _10467_ (.A(_04648_),
    .X(_04649_));
 sky130_fd_sc_hd__mux2_1 _10468_ (.A0(_04636_),
    .A1(_04647_),
    .S(_04649_),
    .X(_04650_));
 sky130_fd_sc_hd__mux2_1 _10469_ (.A0(_01736_),
    .A1(_01898_),
    .S(_01686_),
    .X(_04651_));
 sky130_fd_sc_hd__mux2_1 _10470_ (.A0(_01747_),
    .A1(_01717_),
    .S(_01685_),
    .X(_04652_));
 sky130_fd_sc_hd__mux2_1 _10471_ (.A0(_04651_),
    .A1(_04652_),
    .S(_04628_),
    .X(_04653_));
 sky130_fd_sc_hd__mux2_1 _10472_ (.A0(\leorv32_alu.input1[20] ),
    .A1(_01749_),
    .S(_01685_),
    .X(_04654_));
 sky130_fd_sc_hd__mux2_1 _10473_ (.A0(_01764_),
    .A1(\leorv32_alu.input1[27] ),
    .S(_01685_),
    .X(_04655_));
 sky130_fd_sc_hd__mux2_1 _10474_ (.A0(_04654_),
    .A1(_04655_),
    .S(_04626_),
    .X(_04656_));
 sky130_fd_sc_hd__mux2_1 _10475_ (.A0(_04653_),
    .A1(_04656_),
    .S(_04634_),
    .X(_04657_));
 sky130_fd_sc_hd__mux2_1 _10476_ (.A0(_01868_),
    .A1(_01870_),
    .S(_04624_),
    .X(_04658_));
 sky130_fd_sc_hd__mux2_2 _10477_ (.A0(\leorv32_alu.input1[0] ),
    .A1(\leorv32_alu.input1[31] ),
    .S(\J_type_imm[14] ),
    .X(_04659_));
 sky130_fd_sc_hd__mux2_1 _10478_ (.A0(_04658_),
    .A1(_04659_),
    .S(_04627_),
    .X(_04660_));
 sky130_fd_sc_hd__mux2_1 _10479_ (.A0(\leorv32_alu.input1[24] ),
    .A1(_01784_),
    .S(_01686_),
    .X(_04661_));
 sky130_fd_sc_hd__mux2_1 _10480_ (.A0(\leorv32_alu.input1[8] ),
    .A1(\leorv32_alu.input1[23] ),
    .S(_04624_),
    .X(_04662_));
 sky130_fd_sc_hd__mux2_1 _10481_ (.A0(_04661_),
    .A1(_04662_),
    .S(_04628_),
    .X(_04663_));
 sky130_fd_sc_hd__mux2_1 _10482_ (.A0(_04660_),
    .A1(_04663_),
    .S(_04646_),
    .X(_04664_));
 sky130_fd_sc_hd__clkbuf_4 _10483_ (.A(_04648_),
    .X(_04665_));
 sky130_fd_sc_hd__mux2_1 _10484_ (.A0(_04657_),
    .A1(_04664_),
    .S(_04665_),
    .X(_04666_));
 sky130_fd_sc_hd__or2b_1 _10485_ (.A(_04666_),
    .B_N(_04621_),
    .X(_04667_));
 sky130_fd_sc_hd__o21ai_1 _10486_ (.A1(_04622_),
    .A2(_04650_),
    .B1(_04667_),
    .Y(_04668_));
 sky130_fd_sc_hd__mux2_1 _10487_ (.A0(_01717_),
    .A1(_01747_),
    .S(_01685_),
    .X(_04669_));
 sky130_fd_sc_hd__mux2_1 _10488_ (.A0(_01898_),
    .A1(_01736_),
    .S(\J_type_imm[14] ),
    .X(_04670_));
 sky130_fd_sc_hd__mux2_1 _10489_ (.A0(_04669_),
    .A1(_04670_),
    .S(_04626_),
    .X(_04671_));
 sky130_fd_sc_hd__mux2_1 _10490_ (.A0(\leorv32_alu.input1[27] ),
    .A1(_01764_),
    .S(_01686_),
    .X(_04672_));
 sky130_fd_sc_hd__mux2_1 _10491_ (.A0(_01749_),
    .A1(\leorv32_alu.input1[20] ),
    .S(_01685_),
    .X(_04673_));
 sky130_fd_sc_hd__buf_2 _10492_ (.A(_04626_),
    .X(_04674_));
 sky130_fd_sc_hd__mux2_1 _10493_ (.A0(_04672_),
    .A1(_04673_),
    .S(_04674_),
    .X(_04675_));
 sky130_fd_sc_hd__or2_1 _10494_ (.A(_04635_),
    .B(_04675_),
    .X(_04676_));
 sky130_fd_sc_hd__o21ai_1 _10495_ (.A1(_04646_),
    .A2(_04671_),
    .B1(_04676_),
    .Y(_04677_));
 sky130_fd_sc_hd__mux2_1 _10496_ (.A0(_01711_),
    .A1(_01754_),
    .S(_04624_),
    .X(_04678_));
 sky130_fd_sc_hd__mux2_1 _10497_ (.A0(_01784_),
    .A1(\leorv32_alu.input1[24] ),
    .S(_04624_),
    .X(_04679_));
 sky130_fd_sc_hd__nand2_1 _10498_ (.A(_04674_),
    .B(_04679_),
    .Y(_04680_));
 sky130_fd_sc_hd__o21a_1 _10499_ (.A1(_04674_),
    .A2(_04678_),
    .B1(_04680_),
    .X(_04681_));
 sky130_fd_sc_hd__mux2_1 _10500_ (.A0(\leorv32_alu.input1[31] ),
    .A1(_01807_),
    .S(_01686_),
    .X(_04682_));
 sky130_fd_sc_hd__mux2_1 _10501_ (.A0(_01870_),
    .A1(_01868_),
    .S(_04624_),
    .X(_04683_));
 sky130_fd_sc_hd__mux2_1 _10502_ (.A0(_04682_),
    .A1(_04683_),
    .S(_04628_),
    .X(_04684_));
 sky130_fd_sc_hd__nand2_1 _10503_ (.A(_04646_),
    .B(_04684_),
    .Y(_04685_));
 sky130_fd_sc_hd__inv_2 _10504_ (.A(_04648_),
    .Y(_04686_));
 sky130_fd_sc_hd__clkbuf_4 _10505_ (.A(_04686_),
    .X(_04687_));
 sky130_fd_sc_hd__o211a_1 _10506_ (.A1(_04646_),
    .A2(_04681_),
    .B1(_04685_),
    .C1(_04687_),
    .X(_04688_));
 sky130_fd_sc_hd__a21o_1 _10507_ (.A1(_04649_),
    .A2(_04677_),
    .B1(_04688_),
    .X(_04689_));
 sky130_fd_sc_hd__mux2_1 _10508_ (.A0(_01723_),
    .A1(_01871_),
    .S(\J_type_imm[14] ),
    .X(_04690_));
 sky130_fd_sc_hd__mux2_1 _10509_ (.A0(_01778_),
    .A1(\leorv32_alu.input1[30] ),
    .S(\J_type_imm[14] ),
    .X(_04691_));
 sky130_fd_sc_hd__mux2_1 _10510_ (.A0(_04690_),
    .A1(_04691_),
    .S(_04626_),
    .X(_04692_));
 sky130_fd_sc_hd__mux2_1 _10511_ (.A0(\leorv32_alu.input1[25] ),
    .A1(\leorv32_alu.input1[6] ),
    .S(_01686_),
    .X(_04693_));
 sky130_fd_sc_hd__mux2_1 _10512_ (.A0(_01752_),
    .A1(\leorv32_alu.input1[22] ),
    .S(_01685_),
    .X(_04694_));
 sky130_fd_sc_hd__mux2_1 _10513_ (.A0(_04693_),
    .A1(_04694_),
    .S(_04628_),
    .X(_04695_));
 sky130_fd_sc_hd__or2_1 _10514_ (.A(_04635_),
    .B(_04695_),
    .X(_04696_));
 sky130_fd_sc_hd__o21ai_1 _10515_ (.A1(_04646_),
    .A2(_04692_),
    .B1(_04696_),
    .Y(_04697_));
 sky130_fd_sc_hd__mux2_1 _10516_ (.A0(_01714_),
    .A1(_01880_),
    .S(_04624_),
    .X(_04698_));
 sky130_fd_sc_hd__mux2_1 _10517_ (.A0(\leorv32_alu.input1[5] ),
    .A1(\leorv32_alu.input1[26] ),
    .S(_04624_),
    .X(_04699_));
 sky130_fd_sc_hd__nand2_1 _10518_ (.A(_04674_),
    .B(_04699_),
    .Y(_04700_));
 sky130_fd_sc_hd__o21a_1 _10519_ (.A1(_04674_),
    .A2(_04698_),
    .B1(_04700_),
    .X(_04701_));
 sky130_fd_sc_hd__mux2_1 _10520_ (.A0(\leorv32_alu.input1[29] ),
    .A1(_01901_),
    .S(_01686_),
    .X(_04702_));
 sky130_fd_sc_hd__mux2_1 _10521_ (.A0(_01872_),
    .A1(_01867_),
    .S(_01685_),
    .X(_04703_));
 sky130_fd_sc_hd__mux2_1 _10522_ (.A0(_04702_),
    .A1(_04703_),
    .S(_04628_),
    .X(_04704_));
 sky130_fd_sc_hd__nand2_1 _10523_ (.A(_04646_),
    .B(_04704_),
    .Y(_04705_));
 sky130_fd_sc_hd__o211a_1 _10524_ (.A1(_04646_),
    .A2(_04701_),
    .B1(_04705_),
    .C1(_04687_),
    .X(_04706_));
 sky130_fd_sc_hd__a21o_1 _10525_ (.A1(_04649_),
    .A2(_04697_),
    .B1(_04706_),
    .X(_04707_));
 sky130_fd_sc_hd__clkbuf_4 _10526_ (.A(_04620_),
    .X(_04708_));
 sky130_fd_sc_hd__clkbuf_4 _10527_ (.A(_04708_),
    .X(_04709_));
 sky130_fd_sc_hd__mux2_1 _10528_ (.A0(_04689_),
    .A1(_04707_),
    .S(_04709_),
    .X(_04710_));
 sky130_fd_sc_hd__nand2_2 _10529_ (.A(\barrel_shifter_right.arith ),
    .B(_04659_),
    .Y(_04711_));
 sky130_fd_sc_hd__nand2_2 _10530_ (.A(_04633_),
    .B(_04711_),
    .Y(_04712_));
 sky130_fd_sc_hd__nand2_2 _10531_ (.A(_04626_),
    .B(_04711_),
    .Y(_04713_));
 sky130_fd_sc_hd__buf_2 _10532_ (.A(_04713_),
    .X(_04714_));
 sky130_fd_sc_hd__and3_1 _10533_ (.A(_04659_),
    .B(_04712_),
    .C(_04714_),
    .X(_04715_));
 sky130_fd_sc_hd__nand2_1 _10534_ (.A(_04665_),
    .B(_04711_),
    .Y(_04716_));
 sky130_fd_sc_hd__nand2_1 _10535_ (.A(_04715_),
    .B(_04716_),
    .Y(_04717_));
 sky130_fd_sc_hd__a21o_1 _10536_ (.A1(_04621_),
    .A2(_04711_),
    .B1(_04717_),
    .X(_04718_));
 sky130_fd_sc_hd__clkinv_2 _10537_ (.A(_01564_),
    .Y(_04719_));
 sky130_fd_sc_hd__mux2_1 _10538_ (.A0(_01806_),
    .A1(_04719_),
    .S(_04363_),
    .X(_04720_));
 sky130_fd_sc_hd__buf_2 _10539_ (.A(_04720_),
    .X(_04721_));
 sky130_fd_sc_hd__mux4_1 _10540_ (.A0(_04668_),
    .A1(_04710_),
    .A2(_04711_),
    .A3(_04718_),
    .S0(_04721_),
    .S1(_01688_),
    .X(_04722_));
 sky130_fd_sc_hd__buf_2 _10541_ (.A(_01829_),
    .X(_04723_));
 sky130_fd_sc_hd__nand2_1 _10542_ (.A(_01827_),
    .B(_04420_),
    .Y(_04724_));
 sky130_fd_sc_hd__o211a_1 _10543_ (.A1(_04723_),
    .A2(_04420_),
    .B1(_04724_),
    .C1(_01971_),
    .X(_04725_));
 sky130_fd_sc_hd__o22a_1 _10544_ (.A1(_04619_),
    .A2(_04722_),
    .B1(_04725_),
    .B2(_04419_),
    .X(_04726_));
 sky130_fd_sc_hd__a21o_1 _10545_ (.A1(_04365_),
    .A2(_04617_),
    .B1(_04363_),
    .X(_04727_));
 sky130_fd_sc_hd__nor2_2 _10546_ (.A(_04363_),
    .B(_04365_),
    .Y(_04728_));
 sky130_fd_sc_hd__nor2_4 _10547_ (.A(_04177_),
    .B(_04728_),
    .Y(_04729_));
 sky130_fd_sc_hd__a21oi_1 _10548_ (.A1(_04421_),
    .A2(_04727_),
    .B1(_04729_),
    .Y(_04730_));
 sky130_fd_sc_hd__a31o_1 _10549_ (.A1(_04402_),
    .A2(_04616_),
    .A3(_04726_),
    .B1(_04730_),
    .X(_04731_));
 sky130_fd_sc_hd__a21bo_1 _10550_ (.A1(_04376_),
    .A2(_04400_),
    .B1_N(_04731_),
    .X(_04732_));
 sky130_fd_sc_hd__buf_2 _10551_ (.A(_04182_),
    .X(_04733_));
 sky130_fd_sc_hd__and3_2 _10552_ (.A(_01828_),
    .B(_01903_),
    .C(_04053_),
    .X(_04734_));
 sky130_fd_sc_hd__mux2_1 _10553_ (.A0(net32),
    .A1(net18),
    .S(_04034_),
    .X(_04735_));
 sky130_fd_sc_hd__o21a_2 _10554_ (.A1(_01689_),
    .A2(_04054_),
    .B1(_01970_),
    .X(_04736_));
 sky130_fd_sc_hd__a21oi_1 _10555_ (.A1(_02386_),
    .A2(_04034_),
    .B1(_04736_),
    .Y(_04737_));
 sky130_fd_sc_hd__o21a_1 _10556_ (.A1(net2),
    .A2(_04034_),
    .B1(_04737_),
    .X(_04738_));
 sky130_fd_sc_hd__a221o_1 _10557_ (.A1(net2),
    .A2(_04733_),
    .B1(_04734_),
    .B2(_04735_),
    .C1(_04738_),
    .X(_04739_));
 sky130_fd_sc_hd__and4b_1 _10558_ (.A_N(_01530_),
    .B(\core_state[3] ),
    .C(_01854_),
    .D(_04040_),
    .X(_04740_));
 sky130_fd_sc_hd__buf_2 _10559_ (.A(_04740_),
    .X(_04741_));
 sky130_fd_sc_hd__and2_1 _10560_ (.A(_01527_),
    .B(_04741_),
    .X(_04742_));
 sky130_fd_sc_hd__buf_2 _10561_ (.A(_04742_),
    .X(_04743_));
 sky130_fd_sc_hd__a22o_1 _10562_ (.A1(_04373_),
    .A2(_04732_),
    .B1(_04739_),
    .B2(_04743_),
    .X(_04744_));
 sky130_fd_sc_hd__nand2_1 _10563_ (.A(_01526_),
    .B(_04741_),
    .Y(_04745_));
 sky130_fd_sc_hd__or4_1 _10564_ (.A(_01898_),
    .B(_01901_),
    .C(_01778_),
    .D(_01807_),
    .X(_04746_));
 sky130_fd_sc_hd__or4_1 _10565_ (.A(_01784_),
    .B(\leorv32_alu.input1[6] ),
    .C(\leorv32_alu.input1[5] ),
    .D(_01764_),
    .X(_04747_));
 sky130_fd_sc_hd__or4_1 _10566_ (.A(_01869_),
    .B(_01874_),
    .C(_04746_),
    .D(_04747_),
    .X(_04748_));
 sky130_fd_sc_hd__or4_1 _10567_ (.A(_01749_),
    .B(_01877_),
    .C(_01752_),
    .D(\leorv32_alu.input1[8] ),
    .X(_04749_));
 sky130_fd_sc_hd__or4_1 _10568_ (.A(\leorv32_alu.input1[25] ),
    .B(\leorv32_alu.input1[24] ),
    .C(\leorv32_alu.input1[23] ),
    .D(\leorv32_alu.input1[22] ),
    .X(_04750_));
 sky130_fd_sc_hd__or4_1 _10569_ (.A(\leorv32_alu.input1[29] ),
    .B(_01736_),
    .C(\leorv32_alu.input1[27] ),
    .D(\leorv32_alu.input1[26] ),
    .X(_04751_));
 sky130_fd_sc_hd__or4_1 _10570_ (.A(\leorv32_alu.input1[31] ),
    .B(\leorv32_alu.input1[30] ),
    .C(_01863_),
    .D(_04751_),
    .X(_04752_));
 sky130_fd_sc_hd__or4_2 _10571_ (.A(_04748_),
    .B(_04749_),
    .C(_04750_),
    .D(_04752_),
    .X(_04753_));
 sky130_fd_sc_hd__a41o_1 _10572_ (.A1(\instr[6] ),
    .A2(\instr[5] ),
    .A3(_01530_),
    .A4(_04753_),
    .B1(_04372_),
    .X(_04754_));
 sky130_fd_sc_hd__buf_8 _10573_ (.A(net36),
    .X(_04755_));
 sky130_fd_sc_hd__a21oi_4 _10574_ (.A1(_04745_),
    .A2(_04754_),
    .B1(_04755_),
    .Y(_04756_));
 sky130_fd_sc_hd__or3_4 _10575_ (.A(_02313_),
    .B(_02315_),
    .C(_02241_),
    .X(_04757_));
 sky130_fd_sc_hd__o21a_4 _10576_ (.A1(_01648_),
    .A2(_01642_),
    .B1(_04756_),
    .X(_04758_));
 sky130_fd_sc_hd__a21o_2 _10577_ (.A1(_04756_),
    .A2(_04757_),
    .B1(_04758_),
    .X(_04759_));
 sky130_fd_sc_hd__clkbuf_2 _10578_ (.A(_04759_),
    .X(_04760_));
 sky130_fd_sc_hd__and2_2 _10579_ (.A(_04744_),
    .B(_04760_),
    .X(_04761_));
 sky130_fd_sc_hd__buf_2 _10580_ (.A(_04761_),
    .X(_04762_));
 sky130_fd_sc_hd__nand2_1 _10581_ (.A(_01642_),
    .B(_04756_),
    .Y(_04763_));
 sky130_fd_sc_hd__nor2_2 _10582_ (.A(_01648_),
    .B(_04763_),
    .Y(_04764_));
 sky130_fd_sc_hd__buf_4 _10583_ (.A(_04756_),
    .X(_04765_));
 sky130_fd_sc_hd__nand2_1 _10584_ (.A(_02315_),
    .B(_04765_),
    .Y(_04766_));
 sky130_fd_sc_hd__nor3_4 _10585_ (.A(_02313_),
    .B(_02241_),
    .C(_04766_),
    .Y(_04767_));
 sky130_fd_sc_hd__nand2_4 _10586_ (.A(_04764_),
    .B(_04767_),
    .Y(_04768_));
 sky130_fd_sc_hd__buf_6 _10587_ (.A(_04768_),
    .X(_04769_));
 sky130_fd_sc_hd__mux2_1 _10588_ (.A0(_04762_),
    .A1(\regs[9][0] ),
    .S(_04769_),
    .X(_04770_));
 sky130_fd_sc_hd__clkbuf_1 _10589_ (.A(_04770_),
    .X(_00319_));
 sky130_fd_sc_hd__buf_2 _10590_ (.A(_04759_),
    .X(_04771_));
 sky130_fd_sc_hd__o21ai_4 _10591_ (.A1(_04034_),
    .A2(_04736_),
    .B1(_04173_),
    .Y(_04772_));
 sky130_fd_sc_hd__and2b_1 _10592_ (.A_N(_04736_),
    .B(_04034_),
    .X(_04773_));
 sky130_fd_sc_hd__mux2_1 _10593_ (.A0(net33),
    .A1(net19),
    .S(_04034_),
    .X(_04774_));
 sky130_fd_sc_hd__and2_1 _10594_ (.A(_04734_),
    .B(_04774_),
    .X(_04775_));
 sky130_fd_sc_hd__a221o_1 _10595_ (.A1(net13),
    .A2(_04772_),
    .B1(_04773_),
    .B2(net10),
    .C1(_04775_),
    .X(_04776_));
 sky130_fd_sc_hd__a22o_1 _10596_ (.A1(\instret[1] ),
    .A2(_04384_),
    .B1(_04395_),
    .B2(\instret[33] ),
    .X(_04777_));
 sky130_fd_sc_hd__a221o_1 _10597_ (.A1(\cycles[1] ),
    .A2(_04393_),
    .B1(_04390_),
    .B2(\cycles[33] ),
    .C1(_04777_),
    .X(_04778_));
 sky130_fd_sc_hd__and2_1 _10598_ (.A(_01879_),
    .B(_04617_),
    .X(_04779_));
 sky130_fd_sc_hd__or2_2 _10599_ (.A(_04363_),
    .B(_04779_),
    .X(_04780_));
 sky130_fd_sc_hd__nand2_1 _10600_ (.A(_04366_),
    .B(_04780_),
    .Y(_04781_));
 sky130_fd_sc_hd__buf_4 _10601_ (.A(_04781_),
    .X(_04782_));
 sky130_fd_sc_hd__a21oi_1 _10602_ (.A1(_04417_),
    .A2(_04420_),
    .B1(_04782_),
    .Y(_04783_));
 sky130_fd_sc_hd__o21a_1 _10603_ (.A1(_04417_),
    .A2(_04420_),
    .B1(_04783_),
    .X(_04784_));
 sky130_fd_sc_hd__or4b_1 _10604_ (.A(_01807_),
    .B(_04415_),
    .C(_04416_),
    .D_N(_04418_),
    .X(_04785_));
 sky130_fd_sc_hd__nand2_4 _10605_ (.A(_01602_),
    .B(_04617_),
    .Y(_04786_));
 sky130_fd_sc_hd__nor2_4 _10606_ (.A(_04520_),
    .B(_04786_),
    .Y(_04787_));
 sky130_fd_sc_hd__a31o_1 _10607_ (.A1(_04430_),
    .A2(_04785_),
    .A3(_04787_),
    .B1(_04729_),
    .X(_04788_));
 sky130_fd_sc_hd__nand2_1 _10608_ (.A(_01687_),
    .B(_04617_),
    .Y(_04789_));
 sky130_fd_sc_hd__buf_2 _10609_ (.A(_04789_),
    .X(_04790_));
 sky130_fd_sc_hd__buf_2 _10610_ (.A(_04790_),
    .X(_04791_));
 sky130_fd_sc_hd__o21ai_1 _10611_ (.A1(_04628_),
    .A2(_04683_),
    .B1(_04714_),
    .Y(_04792_));
 sky130_fd_sc_hd__mux2_1 _10612_ (.A0(_04681_),
    .A1(_04792_),
    .S(_04634_),
    .X(_04793_));
 sky130_fd_sc_hd__mux2_1 _10613_ (.A0(_04677_),
    .A1(_04793_),
    .S(_04649_),
    .X(_04794_));
 sky130_fd_sc_hd__mux2_1 _10614_ (.A0(_04707_),
    .A1(_04794_),
    .S(_04621_),
    .X(_04795_));
 sky130_fd_sc_hd__mux2_1 _10615_ (.A0(\rs2_content[0] ),
    .A1(_01564_),
    .S(_04363_),
    .X(_04796_));
 sky130_fd_sc_hd__buf_2 _10616_ (.A(_04796_),
    .X(_04797_));
 sky130_fd_sc_hd__buf_2 _10617_ (.A(_04797_),
    .X(_04798_));
 sky130_fd_sc_hd__mux2_1 _10618_ (.A0(_04668_),
    .A1(_04795_),
    .S(_04798_),
    .X(_04799_));
 sky130_fd_sc_hd__or2_1 _10619_ (.A(_01970_),
    .B(_04799_),
    .X(_04800_));
 sky130_fd_sc_hd__buf_2 _10620_ (.A(_04721_),
    .X(_04801_));
 sky130_fd_sc_hd__o21a_1 _10621_ (.A1(_04674_),
    .A2(_04691_),
    .B1(_04714_),
    .X(_04802_));
 sky130_fd_sc_hd__o21a_1 _10622_ (.A1(_04634_),
    .A2(_04802_),
    .B1(_04712_),
    .X(_04803_));
 sky130_fd_sc_hd__o21ai_1 _10623_ (.A1(_04649_),
    .A2(_04803_),
    .B1(_04716_),
    .Y(_04804_));
 sky130_fd_sc_hd__mux2_1 _10624_ (.A0(_04804_),
    .A1(_04711_),
    .S(_04708_),
    .X(_04805_));
 sky130_fd_sc_hd__a21o_1 _10625_ (.A1(_04797_),
    .A2(_04718_),
    .B1(_01968_),
    .X(_04806_));
 sky130_fd_sc_hd__a21o_1 _10626_ (.A1(_04801_),
    .A2(_04805_),
    .B1(_04806_),
    .X(_04807_));
 sky130_fd_sc_hd__nand3_4 _10627_ (.A(_01687_),
    .B(_01689_),
    .C(_01826_),
    .Y(_04808_));
 sky130_fd_sc_hd__mux2_1 _10628_ (.A0(_01829_),
    .A1(_04808_),
    .S(_04415_),
    .X(_04809_));
 sky130_fd_sc_hd__a21o_1 _10629_ (.A1(_01816_),
    .A2(_04809_),
    .B1(_04416_),
    .X(_04810_));
 sky130_fd_sc_hd__o211a_1 _10630_ (.A1(_02306_),
    .A2(_04807_),
    .B1(_04810_),
    .C1(_04401_),
    .X(_04811_));
 sky130_fd_sc_hd__o21ai_1 _10631_ (.A1(_04791_),
    .A2(_04800_),
    .B1(_04811_),
    .Y(_04812_));
 sky130_fd_sc_hd__o21a_1 _10632_ (.A1(_04784_),
    .A2(_04788_),
    .B1(_04812_),
    .X(_04813_));
 sky130_fd_sc_hd__a221o_1 _10633_ (.A1(\PC[1] ),
    .A2(_04371_),
    .B1(_04376_),
    .B2(_04778_),
    .C1(_04813_),
    .X(_04814_));
 sky130_fd_sc_hd__buf_2 _10634_ (.A(\core_state[1] ),
    .X(_04815_));
 sky130_fd_sc_hd__a22o_1 _10635_ (.A1(_04743_),
    .A2(_04776_),
    .B1(_04814_),
    .B2(_04815_),
    .X(_04816_));
 sky130_fd_sc_hd__and2_2 _10636_ (.A(_04771_),
    .B(_04816_),
    .X(_04817_));
 sky130_fd_sc_hd__buf_2 _10637_ (.A(_04817_),
    .X(_04818_));
 sky130_fd_sc_hd__mux2_1 _10638_ (.A0(_04818_),
    .A1(\regs[9][1] ),
    .S(_04769_),
    .X(_04819_));
 sky130_fd_sc_hd__clkbuf_1 _10639_ (.A(_04819_),
    .X(_00320_));
 sky130_fd_sc_hd__mux2_1 _10640_ (.A0(net3),
    .A1(net20),
    .S(_04034_),
    .X(_04820_));
 sky130_fd_sc_hd__and2_1 _10641_ (.A(_04734_),
    .B(_04820_),
    .X(_04821_));
 sky130_fd_sc_hd__a221o_1 _10642_ (.A1(net24),
    .A2(_04772_),
    .B1(_04773_),
    .B2(net11),
    .C1(_04821_),
    .X(_04822_));
 sky130_fd_sc_hd__a22o_1 _10643_ (.A1(\cycles[34] ),
    .A2(_04390_),
    .B1(_04395_),
    .B2(\instret[34] ),
    .X(_04823_));
 sky130_fd_sc_hd__a221o_1 _10644_ (.A1(\instret[2] ),
    .A2(_04385_),
    .B1(_04393_),
    .B2(\cycles[2] ),
    .C1(_04823_),
    .X(_04824_));
 sky130_fd_sc_hd__clkbuf_4 _10645_ (.A(_04370_),
    .X(_04825_));
 sky130_fd_sc_hd__mux2_1 _10646_ (.A0(_01532_),
    .A1(_04825_),
    .S(_01585_),
    .X(_04826_));
 sky130_fd_sc_hd__clkbuf_4 _10647_ (.A(_04808_),
    .X(_04827_));
 sky130_fd_sc_hd__nor2_1 _10648_ (.A(_01773_),
    .B(_04427_),
    .Y(_04828_));
 sky130_fd_sc_hd__mux2_1 _10649_ (.A0(_04723_),
    .A1(_04827_),
    .S(_04828_),
    .X(_04829_));
 sky130_fd_sc_hd__a22o_1 _10650_ (.A1(_01773_),
    .A2(_04427_),
    .B1(_04829_),
    .B2(_01971_),
    .X(_04830_));
 sky130_fd_sc_hd__clkbuf_4 _10651_ (.A(_01828_),
    .X(_04831_));
 sky130_fd_sc_hd__nor2_1 _10652_ (.A(_02306_),
    .B(_04831_),
    .Y(_04832_));
 sky130_fd_sc_hd__o21a_1 _10653_ (.A1(_04674_),
    .A2(_04638_),
    .B1(_04714_),
    .X(_04833_));
 sky130_fd_sc_hd__o21a_1 _10654_ (.A1(_04635_),
    .A2(_04833_),
    .B1(_04712_),
    .X(_04834_));
 sky130_fd_sc_hd__o21ai_1 _10655_ (.A1(_04649_),
    .A2(_04834_),
    .B1(_04716_),
    .Y(_04835_));
 sky130_fd_sc_hd__mux2_1 _10656_ (.A0(_04835_),
    .A1(_04717_),
    .S(_04708_),
    .X(_04836_));
 sky130_fd_sc_hd__mux2_1 _10657_ (.A0(_04805_),
    .A1(_04836_),
    .S(_04721_),
    .X(_04837_));
 sky130_fd_sc_hd__or2_1 _10658_ (.A(_01969_),
    .B(_04837_),
    .X(_04838_));
 sky130_fd_sc_hd__o21a_1 _10659_ (.A1(_04627_),
    .A2(_04625_),
    .B1(_04713_),
    .X(_04839_));
 sky130_fd_sc_hd__mux2_1 _10660_ (.A0(_04632_),
    .A1(_04839_),
    .S(_04635_),
    .X(_04840_));
 sky130_fd_sc_hd__mux2_1 _10661_ (.A0(_04647_),
    .A1(_04840_),
    .S(_04649_),
    .X(_04841_));
 sky130_fd_sc_hd__mux2_1 _10662_ (.A0(_04666_),
    .A1(_04841_),
    .S(_04709_),
    .X(_04842_));
 sky130_fd_sc_hd__nor2_1 _10663_ (.A(_04801_),
    .B(_04842_),
    .Y(_04843_));
 sky130_fd_sc_hd__a211o_1 _10664_ (.A1(_04801_),
    .A2(_04795_),
    .B1(_04843_),
    .C1(_01969_),
    .X(_04844_));
 sky130_fd_sc_hd__a221o_1 _10665_ (.A1(_04832_),
    .A2(_04838_),
    .B1(_04844_),
    .B2(_02307_),
    .C1(_04618_),
    .X(_04845_));
 sky130_fd_sc_hd__a21o_1 _10666_ (.A1(_04413_),
    .A2(_04414_),
    .B1(_01778_),
    .X(_04846_));
 sky130_fd_sc_hd__a31o_1 _10667_ (.A1(_01807_),
    .A2(_04846_),
    .A3(_04418_),
    .B1(_04415_),
    .X(_04847_));
 sky130_fd_sc_hd__and2_1 _10668_ (.A(_04428_),
    .B(_04847_),
    .X(_04848_));
 sky130_fd_sc_hd__nor2_1 _10669_ (.A(_04428_),
    .B(_04847_),
    .Y(_04849_));
 sky130_fd_sc_hd__or2_2 _10670_ (.A(_04520_),
    .B(_04786_),
    .X(_04850_));
 sky130_fd_sc_hd__a31o_1 _10671_ (.A1(_04428_),
    .A2(_04430_),
    .A3(_04431_),
    .B1(_04850_),
    .X(_04851_));
 sky130_fd_sc_hd__o32a_1 _10672_ (.A1(_04782_),
    .A2(_04848_),
    .A3(_04849_),
    .B1(_04851_),
    .B2(_04432_),
    .X(_04852_));
 sky130_fd_sc_hd__nand2_8 _10673_ (.A(_04401_),
    .B(_04366_),
    .Y(_04853_));
 sky130_fd_sc_hd__a22oi_2 _10674_ (.A1(_04830_),
    .A2(_04845_),
    .B1(_04852_),
    .B2(_04853_),
    .Y(_04854_));
 sky130_fd_sc_hd__a211o_1 _10675_ (.A1(_04376_),
    .A2(_04824_),
    .B1(_04826_),
    .C1(_04854_),
    .X(_04855_));
 sky130_fd_sc_hd__a22o_1 _10676_ (.A1(_04743_),
    .A2(_04822_),
    .B1(_04855_),
    .B2(_04815_),
    .X(_04856_));
 sky130_fd_sc_hd__and2_2 _10677_ (.A(_04771_),
    .B(_04856_),
    .X(_04857_));
 sky130_fd_sc_hd__buf_2 _10678_ (.A(_04857_),
    .X(_04858_));
 sky130_fd_sc_hd__mux2_1 _10679_ (.A0(_04858_),
    .A1(\regs[9][2] ),
    .S(_04769_),
    .X(_04859_));
 sky130_fd_sc_hd__clkbuf_1 _10680_ (.A(_04859_),
    .X(_00321_));
 sky130_fd_sc_hd__mux2_1 _10681_ (.A0(net4),
    .A1(net21),
    .S(_04033_),
    .X(_04860_));
 sky130_fd_sc_hd__and2_1 _10682_ (.A(_04734_),
    .B(_04860_),
    .X(_04861_));
 sky130_fd_sc_hd__a221o_1 _10683_ (.A1(net27),
    .A2(_04772_),
    .B1(_04773_),
    .B2(net12),
    .C1(_04861_),
    .X(_04862_));
 sky130_fd_sc_hd__clkbuf_4 _10684_ (.A(_04825_),
    .X(_04863_));
 sky130_fd_sc_hd__clkbuf_4 _10685_ (.A(_04729_),
    .X(_04864_));
 sky130_fd_sc_hd__o21ai_1 _10686_ (.A1(_04828_),
    .A2(_04848_),
    .B1(_04424_),
    .Y(_04865_));
 sky130_fd_sc_hd__nor2_1 _10687_ (.A(_04363_),
    .B(_04779_),
    .Y(_04866_));
 sky130_fd_sc_hd__nor2_2 _10688_ (.A(_04728_),
    .B(_04866_),
    .Y(_04867_));
 sky130_fd_sc_hd__buf_4 _10689_ (.A(_04867_),
    .X(_04868_));
 sky130_fd_sc_hd__o311a_1 _10690_ (.A1(_04424_),
    .A2(_04828_),
    .A3(_04848_),
    .B1(_04865_),
    .C1(_04868_),
    .X(_04869_));
 sky130_fd_sc_hd__clkbuf_4 _10691_ (.A(_04850_),
    .X(_04870_));
 sky130_fd_sc_hd__a21oi_1 _10692_ (.A1(_04424_),
    .A2(_04433_),
    .B1(_04870_),
    .Y(_04871_));
 sky130_fd_sc_hd__o21a_1 _10693_ (.A1(_04424_),
    .A2(_04433_),
    .B1(_04871_),
    .X(_04872_));
 sky130_fd_sc_hd__o21a_1 _10694_ (.A1(_04674_),
    .A2(_04670_),
    .B1(_04714_),
    .X(_04873_));
 sky130_fd_sc_hd__o21a_1 _10695_ (.A1(_04635_),
    .A2(_04873_),
    .B1(_04712_),
    .X(_04874_));
 sky130_fd_sc_hd__o21ai_1 _10696_ (.A1(_04649_),
    .A2(_04874_),
    .B1(_04716_),
    .Y(_04875_));
 sky130_fd_sc_hd__or2b_1 _10697_ (.A(_04804_),
    .B_N(_04621_),
    .X(_04876_));
 sky130_fd_sc_hd__o21ai_1 _10698_ (.A1(_04709_),
    .A2(_04875_),
    .B1(_04876_),
    .Y(_04877_));
 sky130_fd_sc_hd__nand2_1 _10699_ (.A(_04797_),
    .B(_04836_),
    .Y(_04878_));
 sky130_fd_sc_hd__clkbuf_4 _10700_ (.A(_01817_),
    .X(_04879_));
 sky130_fd_sc_hd__o211a_1 _10701_ (.A1(_04798_),
    .A2(_04877_),
    .B1(_04878_),
    .C1(_04879_),
    .X(_04880_));
 sky130_fd_sc_hd__inv_2 _10702_ (.A(_04880_),
    .Y(_04881_));
 sky130_fd_sc_hd__buf_2 _10703_ (.A(_04797_),
    .X(_04882_));
 sky130_fd_sc_hd__o21a_1 _10704_ (.A1(_04627_),
    .A2(_04703_),
    .B1(_04713_),
    .X(_04883_));
 sky130_fd_sc_hd__clkinv_2 _10705_ (.A(_04883_),
    .Y(_04884_));
 sky130_fd_sc_hd__mux2_1 _10706_ (.A0(_04701_),
    .A1(_04884_),
    .S(_04634_),
    .X(_04885_));
 sky130_fd_sc_hd__mux2_1 _10707_ (.A0(_04697_),
    .A1(_04885_),
    .S(_04649_),
    .X(_04886_));
 sky130_fd_sc_hd__mux2_1 _10708_ (.A0(_04794_),
    .A1(_04886_),
    .S(_04622_),
    .X(_04887_));
 sky130_fd_sc_hd__nor2_1 _10709_ (.A(_04882_),
    .B(_04842_),
    .Y(_04888_));
 sky130_fd_sc_hd__a211o_1 _10710_ (.A1(_04882_),
    .A2(_04887_),
    .B1(_04888_),
    .C1(_01970_),
    .X(_04889_));
 sky130_fd_sc_hd__o21a_1 _10711_ (.A1(_01829_),
    .A2(_04422_),
    .B1(_01816_),
    .X(_04890_));
 sky130_fd_sc_hd__clkbuf_4 _10712_ (.A(_01827_),
    .X(_04891_));
 sky130_fd_sc_hd__nand2_1 _10713_ (.A(_04891_),
    .B(_04422_),
    .Y(_04892_));
 sky130_fd_sc_hd__o211a_1 _10714_ (.A1(_04423_),
    .A2(_04890_),
    .B1(_04892_),
    .C1(_04401_),
    .X(_04893_));
 sky130_fd_sc_hd__o221ai_2 _10715_ (.A1(_02307_),
    .A2(_04881_),
    .B1(_04889_),
    .B2(_04791_),
    .C1(_04893_),
    .Y(_04894_));
 sky130_fd_sc_hd__o31a_1 _10716_ (.A1(_04864_),
    .A2(_04869_),
    .A3(_04872_),
    .B1(_04894_),
    .X(_04895_));
 sky130_fd_sc_hd__clkbuf_4 _10717_ (.A(_04383_),
    .X(_04896_));
 sky130_fd_sc_hd__clkbuf_4 _10718_ (.A(_04394_),
    .X(_04897_));
 sky130_fd_sc_hd__a22o_1 _10719_ (.A1(\cycles[35] ),
    .A2(_04389_),
    .B1(_04897_),
    .B2(\instret[35] ),
    .X(_04898_));
 sky130_fd_sc_hd__a221o_1 _10720_ (.A1(\instret[3] ),
    .A2(_04896_),
    .B1(_04393_),
    .B2(\cycles[3] ),
    .C1(_04898_),
    .X(_04899_));
 sky130_fd_sc_hd__a2bb2o_1 _10721_ (.A1_N(_01858_),
    .A2_N(_02227_),
    .B1(_04375_),
    .B2(_04899_),
    .X(_04900_));
 sky130_fd_sc_hd__a211o_1 _10722_ (.A1(\PC[3] ),
    .A2(_04863_),
    .B1(_04895_),
    .C1(_04900_),
    .X(_04901_));
 sky130_fd_sc_hd__a22o_1 _10723_ (.A1(_04743_),
    .A2(_04862_),
    .B1(_04901_),
    .B2(_04815_),
    .X(_04902_));
 sky130_fd_sc_hd__and2_2 _10724_ (.A(_04771_),
    .B(_04902_),
    .X(_04903_));
 sky130_fd_sc_hd__buf_2 _10725_ (.A(_04903_),
    .X(_04904_));
 sky130_fd_sc_hd__mux2_1 _10726_ (.A0(_04904_),
    .A1(\regs[9][3] ),
    .S(_04769_),
    .X(_04905_));
 sky130_fd_sc_hd__clkbuf_1 _10727_ (.A(_04905_),
    .X(_00322_));
 sky130_fd_sc_hd__mux2_1 _10728_ (.A0(_01900_),
    .A1(_01772_),
    .S(_04365_),
    .X(_04906_));
 sky130_fd_sc_hd__a21o_1 _10729_ (.A1(_01901_),
    .A2(_04906_),
    .B1(_04422_),
    .X(_04907_));
 sky130_fd_sc_hd__or2_1 _10730_ (.A(_01898_),
    .B(_04411_),
    .X(_04908_));
 sky130_fd_sc_hd__a32o_1 _10731_ (.A1(_04424_),
    .A2(_04428_),
    .A3(_04847_),
    .B1(_04907_),
    .B2(_04908_),
    .X(_04909_));
 sky130_fd_sc_hd__and2_1 _10732_ (.A(_04438_),
    .B(_04909_),
    .X(_04910_));
 sky130_fd_sc_hd__nor2_1 _10733_ (.A(_04438_),
    .B(_04909_),
    .Y(_04911_));
 sky130_fd_sc_hd__o32a_1 _10734_ (.A1(_01773_),
    .A2(_04424_),
    .A3(_04906_),
    .B1(_04411_),
    .B2(_01771_),
    .X(_04912_));
 sky130_fd_sc_hd__a211o_1 _10735_ (.A1(_04430_),
    .A2(_04431_),
    .B1(_04424_),
    .C1(_04428_),
    .X(_04913_));
 sky130_fd_sc_hd__a21oi_2 _10736_ (.A1(_04912_),
    .A2(_04913_),
    .B1(_04438_),
    .Y(_04914_));
 sky130_fd_sc_hd__a31o_1 _10737_ (.A1(_04438_),
    .A2(_04912_),
    .A3(_04913_),
    .B1(_04870_),
    .X(_04915_));
 sky130_fd_sc_hd__o32a_1 _10738_ (.A1(_04782_),
    .A2(_04910_),
    .A3(_04911_),
    .B1(_04914_),
    .B2(_04915_),
    .X(_04916_));
 sky130_fd_sc_hd__clkbuf_4 _10739_ (.A(_02307_),
    .X(_04917_));
 sky130_fd_sc_hd__o21a_1 _10740_ (.A1(_04627_),
    .A2(_04655_),
    .B1(_04713_),
    .X(_04918_));
 sky130_fd_sc_hd__o21a_1 _10741_ (.A1(_04635_),
    .A2(_04918_),
    .B1(_04712_),
    .X(_04919_));
 sky130_fd_sc_hd__mux2_1 _10742_ (.A0(_04715_),
    .A1(_04919_),
    .S(_04687_),
    .X(_04920_));
 sky130_fd_sc_hd__nor2_1 _10743_ (.A(_04622_),
    .B(_04920_),
    .Y(_04921_));
 sky130_fd_sc_hd__a21oi_1 _10744_ (.A1(_04622_),
    .A2(_04835_),
    .B1(_04921_),
    .Y(_04922_));
 sky130_fd_sc_hd__o21a_1 _10745_ (.A1(_04721_),
    .A2(_04877_),
    .B1(_04879_),
    .X(_04923_));
 sky130_fd_sc_hd__o21ai_1 _10746_ (.A1(_04882_),
    .A2(_04922_),
    .B1(_04923_),
    .Y(_04924_));
 sky130_fd_sc_hd__and2_1 _10747_ (.A(_01823_),
    .B(_04924_),
    .X(_04925_));
 sky130_fd_sc_hd__buf_2 _10748_ (.A(_04721_),
    .X(_04926_));
 sky130_fd_sc_hd__o21a_1 _10749_ (.A1(_04627_),
    .A2(_04652_),
    .B1(_04713_),
    .X(_04927_));
 sky130_fd_sc_hd__mux2_1 _10750_ (.A0(_04656_),
    .A1(_04927_),
    .S(_04633_),
    .X(_04928_));
 sky130_fd_sc_hd__mux2_1 _10751_ (.A0(_04664_),
    .A1(_04928_),
    .S(_04665_),
    .X(_04929_));
 sky130_fd_sc_hd__mux2_1 _10752_ (.A0(_04841_),
    .A1(_04929_),
    .S(_04621_),
    .X(_04930_));
 sky130_fd_sc_hd__nor2_1 _10753_ (.A(_04926_),
    .B(_04930_),
    .Y(_04931_));
 sky130_fd_sc_hd__a211o_1 _10754_ (.A1(_04926_),
    .A2(_04887_),
    .B1(_04931_),
    .C1(_01970_),
    .X(_04932_));
 sky130_fd_sc_hd__buf_2 _10755_ (.A(_04790_),
    .X(_04933_));
 sky130_fd_sc_hd__mux2_1 _10756_ (.A0(_04723_),
    .A1(_04827_),
    .S(_04436_),
    .X(_04934_));
 sky130_fd_sc_hd__a21o_1 _10757_ (.A1(_01971_),
    .A2(_04934_),
    .B1(_04437_),
    .X(_04935_));
 sky130_fd_sc_hd__o221a_1 _10758_ (.A1(_04917_),
    .A2(_04925_),
    .B1(_04932_),
    .B2(_04933_),
    .C1(_04935_),
    .X(_04936_));
 sky130_fd_sc_hd__a21oi_1 _10759_ (.A1(_04853_),
    .A2(_04916_),
    .B1(_04936_),
    .Y(_04937_));
 sky130_fd_sc_hd__clkbuf_4 _10760_ (.A(_04374_),
    .X(_04938_));
 sky130_fd_sc_hd__clkbuf_4 _10761_ (.A(_04388_),
    .X(_04939_));
 sky130_fd_sc_hd__a22o_1 _10762_ (.A1(\cycles[36] ),
    .A2(_04939_),
    .B1(_04897_),
    .B2(\instret[36] ),
    .X(_04940_));
 sky130_fd_sc_hd__a221o_1 _10763_ (.A1(\instret[4] ),
    .A2(_04896_),
    .B1(_04393_),
    .B2(\cycles[4] ),
    .C1(_04940_),
    .X(_04941_));
 sky130_fd_sc_hd__nor2_1 _10764_ (.A(_01859_),
    .B(_02215_),
    .Y(_04942_));
 sky130_fd_sc_hd__a221o_1 _10765_ (.A1(\PC[4] ),
    .A2(_04825_),
    .B1(_04938_),
    .B2(_04941_),
    .C1(_04942_),
    .X(_04943_));
 sky130_fd_sc_hd__or3_1 _10766_ (.A(_01528_),
    .B(_04937_),
    .C(_04943_),
    .X(_04944_));
 sky130_fd_sc_hd__buf_2 _10767_ (.A(_04741_),
    .X(_04945_));
 sky130_fd_sc_hd__mux2_1 _10768_ (.A0(net5),
    .A1(net22),
    .S(_04034_),
    .X(_04946_));
 sky130_fd_sc_hd__and2_1 _10769_ (.A(_04734_),
    .B(_04946_),
    .X(_04947_));
 sky130_fd_sc_hd__a221o_1 _10770_ (.A1(net28),
    .A2(_04772_),
    .B1(_04773_),
    .B2(_03299_),
    .C1(_04947_),
    .X(_04948_));
 sky130_fd_sc_hd__buf_2 _10771_ (.A(\core_state[1] ),
    .X(_04949_));
 sky130_fd_sc_hd__a21o_1 _10772_ (.A1(_04945_),
    .A2(_04948_),
    .B1(_04949_),
    .X(_04950_));
 sky130_fd_sc_hd__and3_2 _10773_ (.A(_04760_),
    .B(_04944_),
    .C(_04950_),
    .X(_04951_));
 sky130_fd_sc_hd__buf_2 _10774_ (.A(_04951_),
    .X(_04952_));
 sky130_fd_sc_hd__mux2_1 _10775_ (.A0(_04952_),
    .A1(\regs[9][4] ),
    .S(_04769_),
    .X(_04953_));
 sky130_fd_sc_hd__clkbuf_1 _10776_ (.A(_04953_),
    .X(_00323_));
 sky130_fd_sc_hd__mux2_1 _10777_ (.A0(net6),
    .A1(net23),
    .S(_04033_),
    .X(_04954_));
 sky130_fd_sc_hd__and2_1 _10778_ (.A(_04734_),
    .B(_04954_),
    .X(_04955_));
 sky130_fd_sc_hd__a221o_1 _10779_ (.A1(net29),
    .A2(_04772_),
    .B1(_04773_),
    .B2(_03239_),
    .C1(_04955_),
    .X(_04956_));
 sky130_fd_sc_hd__nor2_1 _10780_ (.A(_01765_),
    .B(_04435_),
    .Y(_04957_));
 sky130_fd_sc_hd__nor2_1 _10781_ (.A(_04914_),
    .B(_04957_),
    .Y(_04958_));
 sky130_fd_sc_hd__a21oi_1 _10782_ (.A1(_04612_),
    .A2(_04958_),
    .B1(_04850_),
    .Y(_04959_));
 sky130_fd_sc_hd__o21a_1 _10783_ (.A1(_04612_),
    .A2(_04958_),
    .B1(_04959_),
    .X(_04960_));
 sky130_fd_sc_hd__o21a_1 _10784_ (.A1(_04436_),
    .A2(_04910_),
    .B1(_04612_),
    .X(_04961_));
 sky130_fd_sc_hd__inv_2 _10785_ (.A(_04961_),
    .Y(_04962_));
 sky130_fd_sc_hd__o311a_1 _10786_ (.A1(_04436_),
    .A2(_04612_),
    .A3(_04910_),
    .B1(_04962_),
    .C1(_04868_),
    .X(_04963_));
 sky130_fd_sc_hd__clkinv_2 _10787_ (.A(_04803_),
    .Y(_04964_));
 sky130_fd_sc_hd__o21a_1 _10788_ (.A1(_04674_),
    .A2(_04699_),
    .B1(_04714_),
    .X(_04965_));
 sky130_fd_sc_hd__o21ai_1 _10789_ (.A1(_04635_),
    .A2(_04965_),
    .B1(_04712_),
    .Y(_04966_));
 sky130_fd_sc_hd__mux2_1 _10790_ (.A0(_04964_),
    .A1(_04966_),
    .S(_04687_),
    .X(_04967_));
 sky130_fd_sc_hd__mux2_1 _10791_ (.A0(_04967_),
    .A1(_04875_),
    .S(_04709_),
    .X(_04968_));
 sky130_fd_sc_hd__nor2_1 _10792_ (.A(_04801_),
    .B(_04922_),
    .Y(_04969_));
 sky130_fd_sc_hd__a211o_1 _10793_ (.A1(_04926_),
    .A2(_04968_),
    .B1(_04969_),
    .C1(_01970_),
    .X(_04970_));
 sky130_fd_sc_hd__o21a_1 _10794_ (.A1(_04627_),
    .A2(_04673_),
    .B1(_04713_),
    .X(_04971_));
 sky130_fd_sc_hd__mux2_1 _10795_ (.A0(_04671_),
    .A1(_04971_),
    .S(_04633_),
    .X(_04972_));
 sky130_fd_sc_hd__inv_2 _10796_ (.A(_04972_),
    .Y(_04973_));
 sky130_fd_sc_hd__mux2_1 _10797_ (.A0(_04793_),
    .A1(_04973_),
    .S(_04648_),
    .X(_04974_));
 sky130_fd_sc_hd__and2b_1 _10798_ (.A_N(_04709_),
    .B(_04886_),
    .X(_04975_));
 sky130_fd_sc_hd__a21oi_1 _10799_ (.A1(_04622_),
    .A2(_04974_),
    .B1(_04975_),
    .Y(_04976_));
 sky130_fd_sc_hd__o21a_1 _10800_ (.A1(_04797_),
    .A2(_04930_),
    .B1(_04879_),
    .X(_04977_));
 sky130_fd_sc_hd__o21ai_1 _10801_ (.A1(_04801_),
    .A2(_04976_),
    .B1(_04977_),
    .Y(_04978_));
 sky130_fd_sc_hd__a31o_1 _10802_ (.A1(_01687_),
    .A2(_04441_),
    .A3(_04407_),
    .B1(_01823_),
    .X(_04979_));
 sky130_fd_sc_hd__and2_1 _10803_ (.A(\leorv32_alu.input1[5] ),
    .B(_04406_),
    .X(_04980_));
 sky130_fd_sc_hd__nor2_1 _10804_ (.A(\leorv32_alu.input1[5] ),
    .B(_04406_),
    .Y(_04981_));
 sky130_fd_sc_hd__o2bb2a_1 _10805_ (.A1_N(_01827_),
    .A2_N(_04980_),
    .B1(_04981_),
    .B2(_01816_),
    .X(_04982_));
 sky130_fd_sc_hd__o211a_1 _10806_ (.A1(_04790_),
    .A2(_04978_),
    .B1(_04979_),
    .C1(_04982_),
    .X(_04983_));
 sky130_fd_sc_hd__o21ai_1 _10807_ (.A1(_02307_),
    .A2(_04970_),
    .B1(_04983_),
    .Y(_04984_));
 sky130_fd_sc_hd__o31a_1 _10808_ (.A1(_04729_),
    .A2(_04960_),
    .A3(_04963_),
    .B1(_04984_),
    .X(_04985_));
 sky130_fd_sc_hd__a22o_1 _10809_ (.A1(\cycles[37] ),
    .A2(_04389_),
    .B1(_04897_),
    .B2(\instret[37] ),
    .X(_04986_));
 sky130_fd_sc_hd__a221o_1 _10810_ (.A1(\instret[5] ),
    .A2(_04384_),
    .B1(_04393_),
    .B2(\cycles[5] ),
    .C1(_04986_),
    .X(_04987_));
 sky130_fd_sc_hd__a2bb2o_1 _10811_ (.A1_N(_01858_),
    .A2_N(_02206_),
    .B1(_04375_),
    .B2(_04987_),
    .X(_04988_));
 sky130_fd_sc_hd__a211o_1 _10812_ (.A1(\PC[5] ),
    .A2(_04863_),
    .B1(_04985_),
    .C1(_04988_),
    .X(_04989_));
 sky130_fd_sc_hd__a22o_1 _10813_ (.A1(_04743_),
    .A2(_04956_),
    .B1(_04989_),
    .B2(_04373_),
    .X(_04990_));
 sky130_fd_sc_hd__and2_2 _10814_ (.A(_04771_),
    .B(_04990_),
    .X(_04991_));
 sky130_fd_sc_hd__buf_2 _10815_ (.A(_04991_),
    .X(_04992_));
 sky130_fd_sc_hd__mux2_1 _10816_ (.A0(_04992_),
    .A1(\regs[9][5] ),
    .S(_04769_),
    .X(_04993_));
 sky130_fd_sc_hd__clkbuf_1 _10817_ (.A(_04993_),
    .X(_00324_));
 sky130_fd_sc_hd__mux2_1 _10818_ (.A0(net7),
    .A1(net25),
    .S(_04033_),
    .X(_04994_));
 sky130_fd_sc_hd__and2_1 _10819_ (.A(_04734_),
    .B(_04994_),
    .X(_04995_));
 sky130_fd_sc_hd__a221o_1 _10820_ (.A1(net30),
    .A2(_04772_),
    .B1(_04773_),
    .B2(net16),
    .C1(_04995_),
    .X(_04996_));
 sky130_fd_sc_hd__o21a_1 _10821_ (.A1(_04627_),
    .A2(_04631_),
    .B1(_04713_),
    .X(_04997_));
 sky130_fd_sc_hd__o21a_1 _10822_ (.A1(_04634_),
    .A2(_04997_),
    .B1(_04712_),
    .X(_04998_));
 sky130_fd_sc_hd__mux2_1 _10823_ (.A0(_04834_),
    .A1(_04998_),
    .S(_04687_),
    .X(_04999_));
 sky130_fd_sc_hd__mux2_1 _10824_ (.A0(_04999_),
    .A1(_04920_),
    .S(_04621_),
    .X(_05000_));
 sky130_fd_sc_hd__nor2_1 _10825_ (.A(_04798_),
    .B(_05000_),
    .Y(_05001_));
 sky130_fd_sc_hd__a211o_1 _10826_ (.A1(_04798_),
    .A2(_04968_),
    .B1(_05001_),
    .C1(_01969_),
    .X(_05002_));
 sky130_fd_sc_hd__o21a_1 _10827_ (.A1(_04627_),
    .A2(_04641_),
    .B1(_04714_),
    .X(_05003_));
 sky130_fd_sc_hd__or2_1 _10828_ (.A(_04634_),
    .B(_04639_),
    .X(_05004_));
 sky130_fd_sc_hd__o21ai_1 _10829_ (.A1(_04645_),
    .A2(_05003_),
    .B1(_05004_),
    .Y(_05005_));
 sky130_fd_sc_hd__clkinv_2 _10830_ (.A(_05005_),
    .Y(_05006_));
 sky130_fd_sc_hd__mux2_1 _10831_ (.A0(_04840_),
    .A1(_05006_),
    .S(_04665_),
    .X(_05007_));
 sky130_fd_sc_hd__mux2_1 _10832_ (.A0(_04929_),
    .A1(_05007_),
    .S(_04621_),
    .X(_05008_));
 sky130_fd_sc_hd__o21a_1 _10833_ (.A1(_04721_),
    .A2(_05008_),
    .B1(_04879_),
    .X(_05009_));
 sky130_fd_sc_hd__o21ai_1 _10834_ (.A1(_04882_),
    .A2(_04976_),
    .B1(_05009_),
    .Y(_05010_));
 sky130_fd_sc_hd__and2_1 _10835_ (.A(\leorv32_alu.input1[6] ),
    .B(_04444_),
    .X(_05011_));
 sky130_fd_sc_hd__mux2_1 _10836_ (.A0(_01829_),
    .A1(_04808_),
    .S(_05011_),
    .X(_05012_));
 sky130_fd_sc_hd__a2bb2o_1 _10837_ (.A1_N(\leorv32_alu.input1[6] ),
    .A2_N(_04444_),
    .B1(_05012_),
    .B2(_01816_),
    .X(_05013_));
 sky130_fd_sc_hd__o221a_1 _10838_ (.A1(_02307_),
    .A2(_05002_),
    .B1(_05010_),
    .B2(_04790_),
    .C1(_05013_),
    .X(_05014_));
 sky130_fd_sc_hd__inv_2 _10839_ (.A(_04445_),
    .Y(_05015_));
 sky130_fd_sc_hd__o311ai_4 _10840_ (.A1(_04442_),
    .A2(_04914_),
    .A3(_04957_),
    .B1(_04407_),
    .C1(_05015_),
    .Y(_05016_));
 sky130_fd_sc_hd__or2_1 _10841_ (.A(_04914_),
    .B(_04957_),
    .X(_05017_));
 sky130_fd_sc_hd__a211o_1 _10842_ (.A1(_04407_),
    .A2(_05017_),
    .B1(_05015_),
    .C1(_04442_),
    .X(_05018_));
 sky130_fd_sc_hd__a31o_1 _10843_ (.A1(_04787_),
    .A2(_05016_),
    .A3(_05018_),
    .B1(_04729_),
    .X(_05019_));
 sky130_fd_sc_hd__o21a_1 _10844_ (.A1(_04980_),
    .A2(_04961_),
    .B1(_04445_),
    .X(_05020_));
 sky130_fd_sc_hd__inv_2 _10845_ (.A(_05020_),
    .Y(_05021_));
 sky130_fd_sc_hd__o311a_1 _10846_ (.A1(_04445_),
    .A2(_04980_),
    .A3(_04961_),
    .B1(_05021_),
    .C1(_04868_),
    .X(_05022_));
 sky130_fd_sc_hd__o2bb2a_1 _10847_ (.A1_N(_04402_),
    .A2_N(_05014_),
    .B1(_05019_),
    .B2(_05022_),
    .X(_05023_));
 sky130_fd_sc_hd__a22o_1 _10848_ (.A1(\cycles[6] ),
    .A2(_04392_),
    .B1(_04389_),
    .B2(\cycles[38] ),
    .X(_05024_));
 sky130_fd_sc_hd__a221o_1 _10849_ (.A1(\instret[6] ),
    .A2(_04384_),
    .B1(_04395_),
    .B2(\instret[38] ),
    .C1(_05024_),
    .X(_05025_));
 sky130_fd_sc_hd__a2bb2o_1 _10850_ (.A1_N(_01858_),
    .A2_N(_02191_),
    .B1(_04375_),
    .B2(_05025_),
    .X(_05026_));
 sky130_fd_sc_hd__a211o_1 _10851_ (.A1(_01591_),
    .A2(_04863_),
    .B1(_05023_),
    .C1(_05026_),
    .X(_05027_));
 sky130_fd_sc_hd__a22o_1 _10852_ (.A1(_04743_),
    .A2(_04996_),
    .B1(_05027_),
    .B2(_04373_),
    .X(_05028_));
 sky130_fd_sc_hd__and2_2 _10853_ (.A(_04771_),
    .B(_05028_),
    .X(_05029_));
 sky130_fd_sc_hd__buf_2 _10854_ (.A(_05029_),
    .X(_05030_));
 sky130_fd_sc_hd__mux2_1 _10855_ (.A0(_05030_),
    .A1(\regs[9][6] ),
    .S(_04769_),
    .X(_05031_));
 sky130_fd_sc_hd__clkbuf_1 _10856_ (.A(_05031_),
    .X(_00325_));
 sky130_fd_sc_hd__a21oi_4 _10857_ (.A1(_04765_),
    .A2(_04757_),
    .B1(_04758_),
    .Y(_05032_));
 sky130_fd_sc_hd__buf_2 _10858_ (.A(_04182_),
    .X(_05033_));
 sky130_fd_sc_hd__nand2_1 _10859_ (.A(_03257_),
    .B(_04033_),
    .Y(_05034_));
 sky130_fd_sc_hd__o21a_1 _10860_ (.A1(net31),
    .A2(_04033_),
    .B1(_05034_),
    .X(_05035_));
 sky130_fd_sc_hd__buf_2 _10861_ (.A(_04879_),
    .X(_05036_));
 sky130_fd_sc_hd__mux2_1 _10862_ (.A0(net8),
    .A1(net26),
    .S(_04033_),
    .X(_05037_));
 sky130_fd_sc_hd__nor2_1 _10863_ (.A(_01823_),
    .B(_04054_),
    .Y(_05038_));
 sky130_fd_sc_hd__a22oi_2 _10864_ (.A1(_04734_),
    .A2(_05037_),
    .B1(_05035_),
    .B2(_05038_),
    .Y(_05039_));
 sky130_fd_sc_hd__inv_2 _10865_ (.A(_05039_),
    .Y(_05040_));
 sky130_fd_sc_hd__a221o_1 _10866_ (.A1(net31),
    .A2(_05033_),
    .B1(_05035_),
    .B2(_05036_),
    .C1(_05040_),
    .X(_05041_));
 sky130_fd_sc_hd__nand2_1 _10867_ (.A(\PC[7] ),
    .B(_04863_),
    .Y(_05042_));
 sky130_fd_sc_hd__o21a_1 _10868_ (.A1(_04628_),
    .A2(_04679_),
    .B1(_04714_),
    .X(_05043_));
 sky130_fd_sc_hd__o211a_1 _10869_ (.A1(_04635_),
    .A2(_05043_),
    .B1(_04712_),
    .C1(_04687_),
    .X(_05044_));
 sky130_fd_sc_hd__a21oi_1 _10870_ (.A1(_04649_),
    .A2(_04874_),
    .B1(_05044_),
    .Y(_05045_));
 sky130_fd_sc_hd__mux2_1 _10871_ (.A0(_05045_),
    .A1(_04967_),
    .S(_04709_),
    .X(_05046_));
 sky130_fd_sc_hd__nor2_1 _10872_ (.A(_04801_),
    .B(_05000_),
    .Y(_05047_));
 sky130_fd_sc_hd__a211o_1 _10873_ (.A1(_04926_),
    .A2(_05046_),
    .B1(_05047_),
    .C1(_01970_),
    .X(_05048_));
 sky130_fd_sc_hd__o21a_1 _10874_ (.A1(_04627_),
    .A2(_04694_),
    .B1(_04713_),
    .X(_05049_));
 sky130_fd_sc_hd__mux2_1 _10875_ (.A0(_04692_),
    .A1(_05049_),
    .S(_04633_),
    .X(_05050_));
 sky130_fd_sc_hd__inv_2 _10876_ (.A(_05050_),
    .Y(_05051_));
 sky130_fd_sc_hd__mux2_1 _10877_ (.A0(_04885_),
    .A1(_05051_),
    .S(_04648_),
    .X(_05052_));
 sky130_fd_sc_hd__mux2_1 _10878_ (.A0(_04974_),
    .A1(_05052_),
    .S(_04708_),
    .X(_05053_));
 sky130_fd_sc_hd__nor2_1 _10879_ (.A(_04798_),
    .B(_05008_),
    .Y(_05054_));
 sky130_fd_sc_hd__a211o_1 _10880_ (.A1(_04882_),
    .A2(_05053_),
    .B1(_05054_),
    .C1(_01969_),
    .X(_05055_));
 sky130_fd_sc_hd__and2_1 _10881_ (.A(\J_type_imm[13] ),
    .B(_01815_),
    .X(_05056_));
 sky130_fd_sc_hd__clkbuf_4 _10882_ (.A(_05056_),
    .X(_05057_));
 sky130_fd_sc_hd__or2_1 _10883_ (.A(_01784_),
    .B(_04403_),
    .X(_05058_));
 sky130_fd_sc_hd__and2_1 _10884_ (.A(_01784_),
    .B(_04403_),
    .X(_05059_));
 sky130_fd_sc_hd__a221o_1 _10885_ (.A1(_05057_),
    .A2(_05058_),
    .B1(_05059_),
    .B2(_04891_),
    .C1(_04177_),
    .X(_05060_));
 sky130_fd_sc_hd__a21oi_1 _10886_ (.A1(_04831_),
    .A2(_04443_),
    .B1(_05060_),
    .Y(_05061_));
 sky130_fd_sc_hd__o21a_1 _10887_ (.A1(_04790_),
    .A2(_05055_),
    .B1(_05061_),
    .X(_05062_));
 sky130_fd_sc_hd__o21ai_2 _10888_ (.A1(_04917_),
    .A2(_05048_),
    .B1(_05062_),
    .Y(_05063_));
 sky130_fd_sc_hd__or2_1 _10889_ (.A(_05011_),
    .B(_05020_),
    .X(_05064_));
 sky130_fd_sc_hd__nand2_1 _10890_ (.A(_04443_),
    .B(_05064_),
    .Y(_05065_));
 sky130_fd_sc_hd__o21a_1 _10891_ (.A1(_04443_),
    .A2(_05064_),
    .B1(_04867_),
    .X(_05066_));
 sky130_fd_sc_hd__or2_1 _10892_ (.A(_01767_),
    .B(_04444_),
    .X(_05067_));
 sky130_fd_sc_hd__nand2_1 _10893_ (.A(_05067_),
    .B(_05016_),
    .Y(_05068_));
 sky130_fd_sc_hd__xnor2_1 _10894_ (.A(_04443_),
    .B(_05068_),
    .Y(_05069_));
 sky130_fd_sc_hd__clkbuf_4 _10895_ (.A(_04787_),
    .X(_05070_));
 sky130_fd_sc_hd__a221o_1 _10896_ (.A1(_05065_),
    .A2(_05066_),
    .B1(_05069_),
    .B2(_05070_),
    .C1(_04729_),
    .X(_05071_));
 sky130_fd_sc_hd__clkbuf_4 _10897_ (.A(_04897_),
    .X(_05072_));
 sky130_fd_sc_hd__clkbuf_4 _10898_ (.A(_04392_),
    .X(_05073_));
 sky130_fd_sc_hd__a22o_1 _10899_ (.A1(\cycles[7] ),
    .A2(_05073_),
    .B1(_04390_),
    .B2(\cycles[39] ),
    .X(_05074_));
 sky130_fd_sc_hd__a221o_1 _10900_ (.A1(\instret[7] ),
    .A2(_04385_),
    .B1(_05072_),
    .B2(\instret[39] ),
    .C1(_05074_),
    .X(_05075_));
 sky130_fd_sc_hd__a22oi_1 _10901_ (.A1(_05063_),
    .A2(_05071_),
    .B1(_05075_),
    .B2(_04376_),
    .Y(_05076_));
 sky130_fd_sc_hd__o211a_1 _10902_ (.A1(_01860_),
    .A2(_02183_),
    .B1(_05042_),
    .C1(_05076_),
    .X(_05077_));
 sky130_fd_sc_hd__o2bb2a_1 _10903_ (.A1_N(_04743_),
    .A2_N(_05041_),
    .B1(_05077_),
    .B2(_04372_),
    .X(_05078_));
 sky130_fd_sc_hd__nor2_2 _10904_ (.A(_05032_),
    .B(_05078_),
    .Y(_05079_));
 sky130_fd_sc_hd__buf_2 _10905_ (.A(_05079_),
    .X(_05080_));
 sky130_fd_sc_hd__mux2_1 _10906_ (.A0(_05080_),
    .A1(\regs[9][7] ),
    .S(_04769_),
    .X(_05081_));
 sky130_fd_sc_hd__clkbuf_1 _10907_ (.A(_05081_),
    .X(_00326_));
 sky130_fd_sc_hd__nor2_2 _10908_ (.A(_02306_),
    .B(_05039_),
    .Y(_05082_));
 sky130_fd_sc_hd__a221o_1 _10909_ (.A1(net32),
    .A2(_04733_),
    .B1(_04735_),
    .B2(_05036_),
    .C1(_05082_),
    .X(_05083_));
 sky130_fd_sc_hd__o21a_1 _10910_ (.A1(_04674_),
    .A2(_04662_),
    .B1(_04714_),
    .X(_05084_));
 sky130_fd_sc_hd__and3_1 _10911_ (.A(_04633_),
    .B(_04659_),
    .C(_04714_),
    .X(_05085_));
 sky130_fd_sc_hd__a21o_1 _10912_ (.A1(_04645_),
    .A2(_05084_),
    .B1(_05085_),
    .X(_05086_));
 sky130_fd_sc_hd__mux2_1 _10913_ (.A0(_04919_),
    .A1(_05086_),
    .S(_04687_),
    .X(_05087_));
 sky130_fd_sc_hd__mux2_1 _10914_ (.A0(_05087_),
    .A1(_04999_),
    .S(_04708_),
    .X(_05088_));
 sky130_fd_sc_hd__nor2_1 _10915_ (.A(_04798_),
    .B(_05088_),
    .Y(_05089_));
 sky130_fd_sc_hd__a211o_1 _10916_ (.A1(_04798_),
    .A2(_05046_),
    .B1(_05089_),
    .C1(_01969_),
    .X(_05090_));
 sky130_fd_sc_hd__clkinv_2 _10917_ (.A(_04928_),
    .Y(_05091_));
 sky130_fd_sc_hd__or2_1 _10918_ (.A(_04634_),
    .B(_04660_),
    .X(_05092_));
 sky130_fd_sc_hd__o21ai_1 _10919_ (.A1(_04646_),
    .A2(_05084_),
    .B1(_05092_),
    .Y(_05093_));
 sky130_fd_sc_hd__mux2_1 _10920_ (.A0(_05091_),
    .A1(_05093_),
    .S(_04665_),
    .X(_05094_));
 sky130_fd_sc_hd__nand2_1 _10921_ (.A(_04708_),
    .B(_05094_),
    .Y(_05095_));
 sky130_fd_sc_hd__o21ai_1 _10922_ (.A1(_04621_),
    .A2(_05007_),
    .B1(_05095_),
    .Y(_05096_));
 sky130_fd_sc_hd__mux2_1 _10923_ (.A0(_05053_),
    .A1(_05096_),
    .S(_04797_),
    .X(_05097_));
 sky130_fd_sc_hd__or2_1 _10924_ (.A(_01969_),
    .B(_05097_),
    .X(_05098_));
 sky130_fd_sc_hd__mux2_1 _10925_ (.A0(_01829_),
    .A1(_04808_),
    .S(_04481_),
    .X(_05099_));
 sky130_fd_sc_hd__a21o_1 _10926_ (.A1(_01971_),
    .A2(_05099_),
    .B1(_04482_),
    .X(_05100_));
 sky130_fd_sc_hd__o221a_1 _10927_ (.A1(_02307_),
    .A2(_05090_),
    .B1(_05098_),
    .B2(_04790_),
    .C1(_05100_),
    .X(_05101_));
 sky130_fd_sc_hd__a311o_1 _10928_ (.A1(_04448_),
    .A2(_05067_),
    .A3(_05016_),
    .B1(_04404_),
    .C1(_04483_),
    .X(_05102_));
 sky130_fd_sc_hd__a31o_1 _10929_ (.A1(_04448_),
    .A2(_05067_),
    .A3(_05016_),
    .B1(_04404_),
    .X(_05103_));
 sky130_fd_sc_hd__nand2_1 _10930_ (.A(_04483_),
    .B(_05103_),
    .Y(_05104_));
 sky130_fd_sc_hd__a31o_1 _10931_ (.A1(_04787_),
    .A2(_05102_),
    .A3(_05104_),
    .B1(_04729_),
    .X(_05105_));
 sky130_fd_sc_hd__nor2_1 _10932_ (.A(_04436_),
    .B(_04980_),
    .Y(_05106_));
 sky130_fd_sc_hd__and2_1 _10933_ (.A(_04443_),
    .B(_04445_),
    .X(_05107_));
 sky130_fd_sc_hd__or3b_1 _10934_ (.A(_04981_),
    .B(_05106_),
    .C_N(_05107_),
    .X(_05108_));
 sky130_fd_sc_hd__a21o_1 _10935_ (.A1(_05058_),
    .A2(_05011_),
    .B1(_05059_),
    .X(_05109_));
 sky130_fd_sc_hd__a41oi_2 _10936_ (.A1(_04438_),
    .A2(_04612_),
    .A3(_04909_),
    .A4(_05107_),
    .B1(_05109_),
    .Y(_05110_));
 sky130_fd_sc_hd__a21boi_2 _10937_ (.A1(_05108_),
    .A2(_05110_),
    .B1_N(_04483_),
    .Y(_05111_));
 sky130_fd_sc_hd__a211o_1 _10938_ (.A1(_05058_),
    .A2(_05064_),
    .B1(_05059_),
    .C1(_04483_),
    .X(_05112_));
 sky130_fd_sc_hd__and3b_1 _10939_ (.A_N(_05111_),
    .B(_05112_),
    .C(_04867_),
    .X(_05113_));
 sky130_fd_sc_hd__o2bb2a_1 _10940_ (.A1_N(_04402_),
    .A2_N(_05101_),
    .B1(_05105_),
    .B2(_05113_),
    .X(_05114_));
 sky130_fd_sc_hd__a22o_1 _10941_ (.A1(\cycles[8] ),
    .A2(_04392_),
    .B1(_04939_),
    .B2(\cycles[40] ),
    .X(_05115_));
 sky130_fd_sc_hd__a221o_1 _10942_ (.A1(\instret[8] ),
    .A2(_04896_),
    .B1(_04395_),
    .B2(\instret[40] ),
    .C1(_05115_),
    .X(_05116_));
 sky130_fd_sc_hd__a22o_1 _10943_ (.A1(_01532_),
    .A2(_02162_),
    .B1(_04938_),
    .B2(_05116_),
    .X(_05117_));
 sky130_fd_sc_hd__a211o_1 _10944_ (.A1(\PC[8] ),
    .A2(_04863_),
    .B1(_05114_),
    .C1(_05117_),
    .X(_05118_));
 sky130_fd_sc_hd__a22o_1 _10945_ (.A1(_04743_),
    .A2(_05083_),
    .B1(_05118_),
    .B2(_04373_),
    .X(_05119_));
 sky130_fd_sc_hd__and2_2 _10946_ (.A(_04771_),
    .B(_05119_),
    .X(_05120_));
 sky130_fd_sc_hd__buf_2 _10947_ (.A(_05120_),
    .X(_05121_));
 sky130_fd_sc_hd__mux2_1 _10948_ (.A0(_05121_),
    .A1(\regs[9][8] ),
    .S(_04769_),
    .X(_05122_));
 sky130_fd_sc_hd__clkbuf_1 _10949_ (.A(_05122_),
    .X(_00327_));
 sky130_fd_sc_hd__a221o_1 _10950_ (.A1(net33),
    .A2(_05033_),
    .B1(_04774_),
    .B2(_05036_),
    .C1(_05082_),
    .X(_05123_));
 sky130_fd_sc_hd__o21a_1 _10951_ (.A1(_04481_),
    .A2(_05111_),
    .B1(_04488_),
    .X(_05124_));
 sky130_fd_sc_hd__or3_1 _10952_ (.A(_04481_),
    .B(_04488_),
    .C(_05111_),
    .X(_05125_));
 sky130_fd_sc_hd__or3b_1 _10953_ (.A(_05124_),
    .B(_04782_),
    .C_N(_05125_),
    .X(_05126_));
 sky130_fd_sc_hd__nor2_1 _10954_ (.A(_04486_),
    .B(_04487_),
    .Y(_05127_));
 sky130_fd_sc_hd__o21ai_1 _10955_ (.A1(_01754_),
    .A2(_04480_),
    .B1(_05102_),
    .Y(_05128_));
 sky130_fd_sc_hd__o21ai_1 _10956_ (.A1(_05127_),
    .A2(_05128_),
    .B1(_05070_),
    .Y(_05129_));
 sky130_fd_sc_hd__a21o_1 _10957_ (.A1(_05127_),
    .A2(_05128_),
    .B1(_05129_),
    .X(_05130_));
 sky130_fd_sc_hd__nor2_1 _10958_ (.A(_04645_),
    .B(_05043_),
    .Y(_05131_));
 sky130_fd_sc_hd__a21oi_1 _10959_ (.A1(_04646_),
    .A2(_04792_),
    .B1(_05131_),
    .Y(_05132_));
 sky130_fd_sc_hd__mux2_1 _10960_ (.A0(_04972_),
    .A1(_05132_),
    .S(_04665_),
    .X(_05133_));
 sky130_fd_sc_hd__nand2_1 _10961_ (.A(_04709_),
    .B(_05133_),
    .Y(_05134_));
 sky130_fd_sc_hd__o21ai_1 _10962_ (.A1(_04709_),
    .A2(_05052_),
    .B1(_05134_),
    .Y(_05135_));
 sky130_fd_sc_hd__nor2_1 _10963_ (.A(_04801_),
    .B(_05135_),
    .Y(_05136_));
 sky130_fd_sc_hd__a211o_1 _10964_ (.A1(_04801_),
    .A2(_05096_),
    .B1(_05136_),
    .C1(_01970_),
    .X(_05137_));
 sky130_fd_sc_hd__mux2_1 _10965_ (.A0(_04802_),
    .A1(_05049_),
    .S(_04645_),
    .X(_05138_));
 sky130_fd_sc_hd__inv_2 _10966_ (.A(_05138_),
    .Y(_05139_));
 sky130_fd_sc_hd__mux2_1 _10967_ (.A0(_04966_),
    .A1(_05139_),
    .S(_04687_),
    .X(_05140_));
 sky130_fd_sc_hd__mux2_1 _10968_ (.A0(_05140_),
    .A1(_05045_),
    .S(_04621_),
    .X(_05141_));
 sky130_fd_sc_hd__nor2_1 _10969_ (.A(_04721_),
    .B(_05088_),
    .Y(_05142_));
 sky130_fd_sc_hd__a211o_1 _10970_ (.A1(_04721_),
    .A2(_05141_),
    .B1(_05142_),
    .C1(_01968_),
    .X(_05143_));
 sky130_fd_sc_hd__or2_1 _10971_ (.A(_02306_),
    .B(_05143_),
    .X(_05144_));
 sky130_fd_sc_hd__or2_1 _10972_ (.A(_01752_),
    .B(_04485_),
    .X(_05145_));
 sky130_fd_sc_hd__and2_1 _10973_ (.A(_01752_),
    .B(_04485_),
    .X(_05146_));
 sky130_fd_sc_hd__a221o_1 _10974_ (.A1(_05057_),
    .A2(_05145_),
    .B1(_05146_),
    .B2(_04891_),
    .C1(_04177_),
    .X(_05147_));
 sky130_fd_sc_hd__a21oi_1 _10975_ (.A1(_04831_),
    .A2(_04488_),
    .B1(_05147_),
    .Y(_05148_));
 sky130_fd_sc_hd__o211a_1 _10976_ (.A1(_04791_),
    .A2(_05137_),
    .B1(_05144_),
    .C1(_05148_),
    .X(_05149_));
 sky130_fd_sc_hd__a31o_1 _10977_ (.A1(_04853_),
    .A2(_05126_),
    .A3(_05130_),
    .B1(_05149_),
    .X(_05150_));
 sky130_fd_sc_hd__a22o_1 _10978_ (.A1(\cycles[9] ),
    .A2(_05073_),
    .B1(_04390_),
    .B2(\cycles[41] ),
    .X(_05151_));
 sky130_fd_sc_hd__a221o_1 _10979_ (.A1(\instret[9] ),
    .A2(_04385_),
    .B1(_05072_),
    .B2(\instret[41] ),
    .C1(_05151_),
    .X(_05152_));
 sky130_fd_sc_hd__a22oi_1 _10980_ (.A1(\PC[9] ),
    .A2(_04825_),
    .B1(_04376_),
    .B2(_05152_),
    .Y(_05153_));
 sky130_fd_sc_hd__o211a_1 _10981_ (.A1(_01860_),
    .A2(_02152_),
    .B1(_05150_),
    .C1(_05153_),
    .X(_05154_));
 sky130_fd_sc_hd__o2bb2a_1 _10982_ (.A1_N(_04743_),
    .A2_N(_05123_),
    .B1(_04372_),
    .B2(_05154_),
    .X(_05155_));
 sky130_fd_sc_hd__nor2_2 _10983_ (.A(_05032_),
    .B(_05155_),
    .Y(_05156_));
 sky130_fd_sc_hd__buf_2 _10984_ (.A(_05156_),
    .X(_05157_));
 sky130_fd_sc_hd__mux2_1 _10985_ (.A0(_05157_),
    .A1(\regs[9][9] ),
    .S(_04769_),
    .X(_05158_));
 sky130_fd_sc_hd__clkbuf_1 _10986_ (.A(_05158_),
    .X(_00328_));
 sky130_fd_sc_hd__mux2_1 _10987_ (.A0(_04833_),
    .A1(_05003_),
    .S(_04645_),
    .X(_05159_));
 sky130_fd_sc_hd__mux2_1 _10988_ (.A0(_04998_),
    .A1(_05159_),
    .S(_04686_),
    .X(_05160_));
 sky130_fd_sc_hd__mux2_1 _10989_ (.A0(_05160_),
    .A1(_05087_),
    .S(_04622_),
    .X(_05161_));
 sky130_fd_sc_hd__nor2_1 _10990_ (.A(_04882_),
    .B(_05161_),
    .Y(_05162_));
 sky130_fd_sc_hd__a211o_1 _10991_ (.A1(_04882_),
    .A2(_05141_),
    .B1(_05162_),
    .C1(_01970_),
    .X(_05163_));
 sky130_fd_sc_hd__mux2_1 _10992_ (.A0(_04839_),
    .A1(_04997_),
    .S(_04634_),
    .X(_05164_));
 sky130_fd_sc_hd__inv_2 _10993_ (.A(_05164_),
    .Y(_05165_));
 sky130_fd_sc_hd__mux2_1 _10994_ (.A0(_05005_),
    .A1(_05165_),
    .S(_04665_),
    .X(_05166_));
 sky130_fd_sc_hd__mux2_1 _10995_ (.A0(_05094_),
    .A1(_05166_),
    .S(_04709_),
    .X(_05167_));
 sky130_fd_sc_hd__nor2_1 _10996_ (.A(_04797_),
    .B(_05135_),
    .Y(_05168_));
 sky130_fd_sc_hd__a211o_1 _10997_ (.A1(_04798_),
    .A2(_05167_),
    .B1(_05168_),
    .C1(_01969_),
    .X(_05169_));
 sky130_fd_sc_hd__mux2_1 _10998_ (.A0(_04723_),
    .A1(_04827_),
    .S(_04471_),
    .X(_05170_));
 sky130_fd_sc_hd__a21o_1 _10999_ (.A1(_01971_),
    .A2(_05170_),
    .B1(_04473_),
    .X(_05171_));
 sky130_fd_sc_hd__o221a_1 _11000_ (.A1(_04917_),
    .A2(_05163_),
    .B1(_05169_),
    .B2(_04791_),
    .C1(_05171_),
    .X(_05172_));
 sky130_fd_sc_hd__o21a_1 _11001_ (.A1(_05146_),
    .A2(_05124_),
    .B1(_04474_),
    .X(_05173_));
 sky130_fd_sc_hd__o31ai_1 _11002_ (.A1(_04474_),
    .A2(_05146_),
    .A3(_05124_),
    .B1(_04868_),
    .Y(_05174_));
 sky130_fd_sc_hd__o22a_1 _11003_ (.A1(_04484_),
    .A2(_04485_),
    .B1(_04480_),
    .B2(_01754_),
    .X(_05175_));
 sky130_fd_sc_hd__a21o_1 _11004_ (.A1(_05102_),
    .A2(_05175_),
    .B1(_04486_),
    .X(_05176_));
 sky130_fd_sc_hd__xor2_1 _11005_ (.A(_04474_),
    .B(_05176_),
    .X(_05177_));
 sky130_fd_sc_hd__a2bb2o_1 _11006_ (.A1_N(_05173_),
    .A2_N(_05174_),
    .B1(_05177_),
    .B2(_05070_),
    .X(_05178_));
 sky130_fd_sc_hd__o2bb2a_1 _11007_ (.A1_N(_04402_),
    .A2_N(_05172_),
    .B1(_04864_),
    .B2(_05178_),
    .X(_05179_));
 sky130_fd_sc_hd__a22o_1 _11008_ (.A1(\cycles[42] ),
    .A2(_04939_),
    .B1(_04897_),
    .B2(\instret[42] ),
    .X(_05180_));
 sky130_fd_sc_hd__a221o_1 _11009_ (.A1(\instret[10] ),
    .A2(_04385_),
    .B1(_04393_),
    .B2(\cycles[10] ),
    .C1(_05180_),
    .X(_05181_));
 sky130_fd_sc_hd__a221o_1 _11010_ (.A1(\PC[10] ),
    .A2(_04863_),
    .B1(_04376_),
    .B2(_05181_),
    .C1(_01527_),
    .X(_05182_));
 sky130_fd_sc_hd__a211o_1 _11011_ (.A1(_01532_),
    .A2(_02140_),
    .B1(_05179_),
    .C1(_05182_),
    .X(_05183_));
 sky130_fd_sc_hd__a221o_1 _11012_ (.A1(net3),
    .A2(_04733_),
    .B1(_04820_),
    .B2(_05036_),
    .C1(_05082_),
    .X(_05184_));
 sky130_fd_sc_hd__a21o_1 _11013_ (.A1(_04945_),
    .A2(_05184_),
    .B1(_04949_),
    .X(_05185_));
 sky130_fd_sc_hd__and3_2 _11014_ (.A(_04760_),
    .B(_05183_),
    .C(_05185_),
    .X(_05186_));
 sky130_fd_sc_hd__clkbuf_4 _11015_ (.A(_05186_),
    .X(_05187_));
 sky130_fd_sc_hd__buf_4 _11016_ (.A(_04768_),
    .X(_05188_));
 sky130_fd_sc_hd__mux2_1 _11017_ (.A0(_05187_),
    .A1(\regs[9][10] ),
    .S(_05188_),
    .X(_05189_));
 sky130_fd_sc_hd__clkbuf_1 _11018_ (.A(_05189_),
    .X(_00329_));
 sky130_fd_sc_hd__nor2_1 _11019_ (.A(_04474_),
    .B(_05176_),
    .Y(_05190_));
 sky130_fd_sc_hd__a21o_1 _11020_ (.A1(_01877_),
    .A2(_04470_),
    .B1(_05190_),
    .X(_05191_));
 sky130_fd_sc_hd__xnor2_1 _11021_ (.A(_04478_),
    .B(_05191_),
    .Y(_05192_));
 sky130_fd_sc_hd__or3_1 _11022_ (.A(_04471_),
    .B(_04478_),
    .C(_05173_),
    .X(_05193_));
 sky130_fd_sc_hd__o21ai_1 _11023_ (.A1(_04471_),
    .A2(_05173_),
    .B1(_04478_),
    .Y(_05194_));
 sky130_fd_sc_hd__and3_1 _11024_ (.A(_04868_),
    .B(_05193_),
    .C(_05194_),
    .X(_05195_));
 sky130_fd_sc_hd__a211o_1 _11025_ (.A1(_05070_),
    .A2(_05192_),
    .B1(_05195_),
    .C1(_04864_),
    .X(_05196_));
 sky130_fd_sc_hd__mux2_1 _11026_ (.A0(_04883_),
    .A1(_04965_),
    .S(_04634_),
    .X(_05197_));
 sky130_fd_sc_hd__mux2_1 _11027_ (.A0(_05050_),
    .A1(_05197_),
    .S(_04665_),
    .X(_05198_));
 sky130_fd_sc_hd__mux2_1 _11028_ (.A0(_05133_),
    .A1(_05198_),
    .S(_04708_),
    .X(_05199_));
 sky130_fd_sc_hd__nor2_1 _11029_ (.A(_04926_),
    .B(_05199_),
    .Y(_05200_));
 sky130_fd_sc_hd__a211o_1 _11030_ (.A1(_04926_),
    .A2(_05167_),
    .B1(_05200_),
    .C1(_01970_),
    .X(_05201_));
 sky130_fd_sc_hd__mux2_1 _11031_ (.A0(_04873_),
    .A1(_04971_),
    .S(_04645_),
    .X(_05202_));
 sky130_fd_sc_hd__o211a_1 _11032_ (.A1(_04635_),
    .A2(_05043_),
    .B1(_04712_),
    .C1(_04648_),
    .X(_05203_));
 sky130_fd_sc_hd__a21o_1 _11033_ (.A1(_04687_),
    .A2(_05202_),
    .B1(_05203_),
    .X(_05204_));
 sky130_fd_sc_hd__nor2_1 _11034_ (.A(_04709_),
    .B(_05204_),
    .Y(_05205_));
 sky130_fd_sc_hd__a21oi_1 _11035_ (.A1(_04622_),
    .A2(_05140_),
    .B1(_05205_),
    .Y(_05206_));
 sky130_fd_sc_hd__o21a_1 _11036_ (.A1(_04926_),
    .A2(_05161_),
    .B1(_04879_),
    .X(_05207_));
 sky130_fd_sc_hd__o21ai_1 _11037_ (.A1(_04882_),
    .A2(_05206_),
    .B1(_05207_),
    .Y(_05208_));
 sky130_fd_sc_hd__o21a_1 _11038_ (.A1(\rs2_content[11] ),
    .A2(_04503_),
    .B1(_04497_),
    .X(_05209_));
 sky130_fd_sc_hd__or2_1 _11039_ (.A(_01749_),
    .B(_05209_),
    .X(_05210_));
 sky130_fd_sc_hd__and2_1 _11040_ (.A(_01749_),
    .B(_05209_),
    .X(_05211_));
 sky130_fd_sc_hd__a221o_1 _11041_ (.A1(_05057_),
    .A2(_05210_),
    .B1(_05211_),
    .B2(_04891_),
    .C1(_04177_),
    .X(_05212_));
 sky130_fd_sc_hd__a21o_1 _11042_ (.A1(_04831_),
    .A2(_04478_),
    .B1(_05212_),
    .X(_05213_));
 sky130_fd_sc_hd__o21ba_1 _11043_ (.A1(_02308_),
    .A2(_05208_),
    .B1_N(_05213_),
    .X(_05214_));
 sky130_fd_sc_hd__o21ai_1 _11044_ (.A1(_04933_),
    .A2(_05201_),
    .B1(_05214_),
    .Y(_05215_));
 sky130_fd_sc_hd__a22o_1 _11045_ (.A1(\cycles[11] ),
    .A2(_05073_),
    .B1(_04939_),
    .B2(\cycles[43] ),
    .X(_05216_));
 sky130_fd_sc_hd__a221o_1 _11046_ (.A1(\instret[11] ),
    .A2(_04896_),
    .B1(_05072_),
    .B2(\instret[43] ),
    .C1(_05216_),
    .X(_05217_));
 sky130_fd_sc_hd__nor2_1 _11047_ (.A(_01859_),
    .B(_02129_),
    .Y(_05218_));
 sky130_fd_sc_hd__a221o_1 _11048_ (.A1(\PC[11] ),
    .A2(_04825_),
    .B1(_04938_),
    .B2(_05217_),
    .C1(_05218_),
    .X(_05219_));
 sky130_fd_sc_hd__a211o_1 _11049_ (.A1(_05196_),
    .A2(_05215_),
    .B1(_05219_),
    .C1(_01528_),
    .X(_05220_));
 sky130_fd_sc_hd__a221o_1 _11050_ (.A1(net4),
    .A2(_04733_),
    .B1(_04860_),
    .B2(_05036_),
    .C1(_05082_),
    .X(_05221_));
 sky130_fd_sc_hd__a21o_1 _11051_ (.A1(_04945_),
    .A2(_05221_),
    .B1(_04949_),
    .X(_05222_));
 sky130_fd_sc_hd__and3_4 _11052_ (.A(_04760_),
    .B(_05220_),
    .C(_05222_),
    .X(_05223_));
 sky130_fd_sc_hd__clkbuf_4 _11053_ (.A(_05223_),
    .X(_05224_));
 sky130_fd_sc_hd__mux2_1 _11054_ (.A0(_05224_),
    .A1(\regs[9][11] ),
    .S(_05188_),
    .X(_05225_));
 sky130_fd_sc_hd__clkbuf_1 _11055_ (.A(_05225_),
    .X(_00330_));
 sky130_fd_sc_hd__a221o_1 _11056_ (.A1(net5),
    .A2(_04733_),
    .B1(_04946_),
    .B2(_05036_),
    .C1(_05082_),
    .X(_05226_));
 sky130_fd_sc_hd__buf_2 _11057_ (.A(_04361_),
    .X(_05227_));
 sky130_fd_sc_hd__a22o_1 _11058_ (.A1(\cycles[44] ),
    .A2(_04388_),
    .B1(_04394_),
    .B2(\instret[44] ),
    .X(_05228_));
 sky130_fd_sc_hd__a221o_1 _11059_ (.A1(\instret[12] ),
    .A2(_04383_),
    .B1(_04392_),
    .B2(\cycles[12] ),
    .C1(_05228_),
    .X(_05229_));
 sky130_fd_sc_hd__and2b_1 _11060_ (.A_N(_02115_),
    .B(_04370_),
    .X(_05230_));
 sky130_fd_sc_hd__a221o_1 _11061_ (.A1(_01826_),
    .A2(_05227_),
    .B1(_04374_),
    .B2(_05229_),
    .C1(_05230_),
    .X(_05231_));
 sky130_fd_sc_hd__nor2_1 _11062_ (.A(_01859_),
    .B(_02083_),
    .Y(_05232_));
 sky130_fd_sc_hd__mux2_1 _11063_ (.A0(_04918_),
    .A1(_04927_),
    .S(_04645_),
    .X(_05233_));
 sky130_fd_sc_hd__clkinv_2 _11064_ (.A(_05233_),
    .Y(_05234_));
 sky130_fd_sc_hd__mux2_1 _11065_ (.A0(_05093_),
    .A1(_05234_),
    .S(_04665_),
    .X(_05235_));
 sky130_fd_sc_hd__mux2_1 _11066_ (.A0(_05166_),
    .A1(_05235_),
    .S(_04708_),
    .X(_05236_));
 sky130_fd_sc_hd__nor2_1 _11067_ (.A(_04797_),
    .B(_05199_),
    .Y(_05237_));
 sky130_fd_sc_hd__a211o_1 _11068_ (.A1(_04798_),
    .A2(_05236_),
    .B1(_05237_),
    .C1(_01969_),
    .X(_05238_));
 sky130_fd_sc_hd__mux2_1 _11069_ (.A0(_05086_),
    .A1(_05233_),
    .S(_04686_),
    .X(_05239_));
 sky130_fd_sc_hd__mux2_1 _11070_ (.A0(_05239_),
    .A1(_05160_),
    .S(_04620_),
    .X(_05240_));
 sky130_fd_sc_hd__o21a_1 _11071_ (.A1(_04797_),
    .A2(_05240_),
    .B1(_04879_),
    .X(_05241_));
 sky130_fd_sc_hd__o21ai_1 _11072_ (.A1(_04801_),
    .A2(_05206_),
    .B1(_05241_),
    .Y(_05242_));
 sky130_fd_sc_hd__mux2_1 _11073_ (.A0(_01829_),
    .A1(_04808_),
    .S(_04465_),
    .X(_05243_));
 sky130_fd_sc_hd__a21o_1 _11074_ (.A1(_01816_),
    .A2(_05243_),
    .B1(_04467_),
    .X(_05244_));
 sky130_fd_sc_hd__o221a_1 _11075_ (.A1(_04790_),
    .A2(_05238_),
    .B1(_05242_),
    .B2(_02306_),
    .C1(_05244_),
    .X(_05245_));
 sky130_fd_sc_hd__and2_1 _11076_ (.A(_04474_),
    .B(_04478_),
    .X(_05246_));
 sky130_fd_sc_hd__o21a_1 _11077_ (.A1(_04481_),
    .A2(_05146_),
    .B1(_05145_),
    .X(_05247_));
 sky130_fd_sc_hd__a221o_1 _11078_ (.A1(_04471_),
    .A2(_05210_),
    .B1(_05246_),
    .B2(_05247_),
    .C1(_05211_),
    .X(_05248_));
 sky130_fd_sc_hd__a31oi_2 _11079_ (.A1(_04488_),
    .A2(_05111_),
    .A3(_05246_),
    .B1(_05248_),
    .Y(_05249_));
 sky130_fd_sc_hd__and2_1 _11080_ (.A(_04468_),
    .B(_05249_),
    .X(_05250_));
 sky130_fd_sc_hd__nor2_1 _11081_ (.A(_04468_),
    .B(_05249_),
    .Y(_05251_));
 sky130_fd_sc_hd__or2_1 _11082_ (.A(_05250_),
    .B(_05251_),
    .X(_05252_));
 sky130_fd_sc_hd__a21o_1 _11083_ (.A1(_01877_),
    .A2(_04470_),
    .B1(_04476_),
    .X(_05253_));
 sky130_fd_sc_hd__o211a_1 _11084_ (.A1(_05190_),
    .A2(_05253_),
    .B1(_04468_),
    .C1(_04477_),
    .X(_05254_));
 sky130_fd_sc_hd__a21o_1 _11085_ (.A1(_04520_),
    .A2(_05252_),
    .B1(_04786_),
    .X(_05255_));
 sky130_fd_sc_hd__a211o_1 _11086_ (.A1(_04477_),
    .A2(_05191_),
    .B1(_04468_),
    .C1(_04476_),
    .X(_05256_));
 sky130_fd_sc_hd__or3b_1 _11087_ (.A(_05254_),
    .B(_05255_),
    .C_N(_05256_),
    .X(_05257_));
 sky130_fd_sc_hd__o211a_1 _11088_ (.A1(_04866_),
    .A2(_05252_),
    .B1(_05257_),
    .C1(_04177_),
    .X(_05258_));
 sky130_fd_sc_hd__a211o_1 _11089_ (.A1(_04401_),
    .A2(_05245_),
    .B1(_05258_),
    .C1(_04728_),
    .X(_05259_));
 sky130_fd_sc_hd__or3b_1 _11090_ (.A(_05231_),
    .B(_05232_),
    .C_N(_05259_),
    .X(_05260_));
 sky130_fd_sc_hd__a22o_1 _11091_ (.A1(_04743_),
    .A2(_05226_),
    .B1(_05260_),
    .B2(_04815_),
    .X(_05261_));
 sky130_fd_sc_hd__and2_4 _11092_ (.A(_04771_),
    .B(_05261_),
    .X(_05262_));
 sky130_fd_sc_hd__buf_2 _11093_ (.A(_05262_),
    .X(_05263_));
 sky130_fd_sc_hd__mux2_1 _11094_ (.A0(_05263_),
    .A1(\regs[9][12] ),
    .S(_05188_),
    .X(_05264_));
 sky130_fd_sc_hd__clkbuf_1 _11095_ (.A(_05264_),
    .X(_00331_));
 sky130_fd_sc_hd__a221o_1 _11096_ (.A1(net6),
    .A2(_04182_),
    .B1(_04954_),
    .B2(_05036_),
    .C1(_05082_),
    .X(_05265_));
 sky130_fd_sc_hd__o21ai_1 _11097_ (.A1(_04465_),
    .A2(_05251_),
    .B1(_04464_),
    .Y(_05266_));
 sky130_fd_sc_hd__or3_1 _11098_ (.A(_04464_),
    .B(_04465_),
    .C(_05251_),
    .X(_05267_));
 sky130_fd_sc_hd__a31o_1 _11099_ (.A1(_04867_),
    .A2(_05266_),
    .A3(_05267_),
    .B1(_04729_),
    .X(_05268_));
 sky130_fd_sc_hd__a21oi_1 _11100_ (.A1(_01747_),
    .A2(_04466_),
    .B1(_05254_),
    .Y(_05269_));
 sky130_fd_sc_hd__o21ai_1 _11101_ (.A1(_04464_),
    .A2(_05269_),
    .B1(_04787_),
    .Y(_05270_));
 sky130_fd_sc_hd__a21oi_1 _11102_ (.A1(_04464_),
    .A2(_05269_),
    .B1(_05270_),
    .Y(_05271_));
 sky130_fd_sc_hd__nor2_1 _11103_ (.A(_01872_),
    .B(_04461_),
    .Y(_05272_));
 sky130_fd_sc_hd__mux2_1 _11104_ (.A0(_05132_),
    .A1(_05202_),
    .S(_04665_),
    .X(_05273_));
 sky130_fd_sc_hd__mux2_1 _11105_ (.A0(_05198_),
    .A1(_05273_),
    .S(_04708_),
    .X(_05274_));
 sky130_fd_sc_hd__nor2_1 _11106_ (.A(_04720_),
    .B(_05274_),
    .Y(_05275_));
 sky130_fd_sc_hd__a211o_1 _11107_ (.A1(_04721_),
    .A2(_05236_),
    .B1(_05275_),
    .C1(_01968_),
    .X(_05276_));
 sky130_fd_sc_hd__nor2_1 _11108_ (.A(_01688_),
    .B(_01823_),
    .Y(_05277_));
 sky130_fd_sc_hd__nand2_1 _11109_ (.A(_05277_),
    .B(_04464_),
    .Y(_05278_));
 sky130_fd_sc_hd__o221ai_1 _11110_ (.A1(_01971_),
    .A2(_05272_),
    .B1(_04790_),
    .B2(_05276_),
    .C1(_05278_),
    .Y(_05279_));
 sky130_fd_sc_hd__nand2_1 _11111_ (.A(_01872_),
    .B(_04461_),
    .Y(_05280_));
 sky130_fd_sc_hd__mux2_1 _11112_ (.A0(_05138_),
    .A1(_05197_),
    .S(_04687_),
    .X(_05281_));
 sky130_fd_sc_hd__mux2_1 _11113_ (.A0(_05281_),
    .A1(_05204_),
    .S(_04708_),
    .X(_05282_));
 sky130_fd_sc_hd__o21a_1 _11114_ (.A1(_04720_),
    .A2(_05240_),
    .B1(_01817_),
    .X(_05283_));
 sky130_fd_sc_hd__o21ai_1 _11115_ (.A1(_04797_),
    .A2(_05282_),
    .B1(_05283_),
    .Y(_05284_));
 sky130_fd_sc_hd__o221a_1 _11116_ (.A1(_04808_),
    .A2(_05280_),
    .B1(_05284_),
    .B2(_01687_),
    .C1(_04401_),
    .X(_05285_));
 sky130_fd_sc_hd__and2b_1 _11117_ (.A_N(_05279_),
    .B(_05285_),
    .X(_05286_));
 sky130_fd_sc_hd__o21ba_1 _11118_ (.A1(_05268_),
    .A2(_05271_),
    .B1_N(_05286_),
    .X(_05287_));
 sky130_fd_sc_hd__a22o_1 _11119_ (.A1(\cycles[13] ),
    .A2(_04391_),
    .B1(_04388_),
    .B2(\cycles[45] ),
    .X(_05288_));
 sky130_fd_sc_hd__a221o_1 _11120_ (.A1(\instret[13] ),
    .A2(_04383_),
    .B1(_04394_),
    .B2(\instret[45] ),
    .C1(_05288_),
    .X(_05289_));
 sky130_fd_sc_hd__a22o_1 _11121_ (.A1(_01689_),
    .A2(_04361_),
    .B1(_04374_),
    .B2(_05289_),
    .X(_05290_));
 sky130_fd_sc_hd__a31o_1 _11122_ (.A1(_01562_),
    .A2(_02107_),
    .A3(_04825_),
    .B1(_05290_),
    .X(_05291_));
 sky130_fd_sc_hd__nor2_1 _11123_ (.A(_01859_),
    .B(_02110_),
    .Y(_05292_));
 sky130_fd_sc_hd__or3_1 _11124_ (.A(_05287_),
    .B(_05291_),
    .C(_05292_),
    .X(_05293_));
 sky130_fd_sc_hd__a22o_1 _11125_ (.A1(_04742_),
    .A2(_05265_),
    .B1(_05293_),
    .B2(_04815_),
    .X(_05294_));
 sky130_fd_sc_hd__and2_2 _11126_ (.A(_04760_),
    .B(_05294_),
    .X(_05295_));
 sky130_fd_sc_hd__clkbuf_4 _11127_ (.A(_05295_),
    .X(_05296_));
 sky130_fd_sc_hd__mux2_1 _11128_ (.A0(_05296_),
    .A1(\regs[9][13] ),
    .S(_05188_),
    .X(_05297_));
 sky130_fd_sc_hd__clkbuf_1 _11129_ (.A(_05297_),
    .X(_00332_));
 sky130_fd_sc_hd__a221o_1 _11130_ (.A1(net7),
    .A2(_04182_),
    .B1(_04994_),
    .B2(_05036_),
    .C1(_05082_),
    .X(_05298_));
 sky130_fd_sc_hd__buf_2 _11131_ (.A(_04825_),
    .X(_05299_));
 sky130_fd_sc_hd__xor2_1 _11132_ (.A(_01614_),
    .B(_02098_),
    .X(_05300_));
 sky130_fd_sc_hd__a22o_1 _11133_ (.A1(\cycles[46] ),
    .A2(_04389_),
    .B1(_04394_),
    .B2(\instret[46] ),
    .X(_05301_));
 sky130_fd_sc_hd__a221o_1 _11134_ (.A1(\instret[14] ),
    .A2(_04384_),
    .B1(_05073_),
    .B2(\cycles[14] ),
    .C1(_05301_),
    .X(_05302_));
 sky130_fd_sc_hd__nor2_1 _11135_ (.A(_01858_),
    .B(_02089_),
    .Y(_05303_));
 sky130_fd_sc_hd__a221o_1 _11136_ (.A1(_04917_),
    .A2(_05227_),
    .B1(_04375_),
    .B2(_05302_),
    .C1(_05303_),
    .X(_05304_));
 sky130_fd_sc_hd__mux2_1 _11137_ (.A0(_05159_),
    .A1(_05164_),
    .S(_04686_),
    .X(_05305_));
 sky130_fd_sc_hd__mux2_1 _11138_ (.A0(_05305_),
    .A1(_05239_),
    .S(_04620_),
    .X(_05306_));
 sky130_fd_sc_hd__o21a_1 _11139_ (.A1(_04796_),
    .A2(_05306_),
    .B1(_01817_),
    .X(_05307_));
 sky130_fd_sc_hd__o21ai_1 _11140_ (.A1(_04721_),
    .A2(_05282_),
    .B1(_05307_),
    .Y(_05308_));
 sky130_fd_sc_hd__nand2_1 _11141_ (.A(_04622_),
    .B(_05305_),
    .Y(_05309_));
 sky130_fd_sc_hd__o21ai_1 _11142_ (.A1(_04622_),
    .A2(_05235_),
    .B1(_05309_),
    .Y(_05310_));
 sky130_fd_sc_hd__o21a_1 _11143_ (.A1(_04798_),
    .A2(_05274_),
    .B1(_04879_),
    .X(_05311_));
 sky130_fd_sc_hd__o21ai_1 _11144_ (.A1(_04801_),
    .A2(_05310_),
    .B1(_05311_),
    .Y(_05312_));
 sky130_fd_sc_hd__mux2_1 _11145_ (.A0(_01829_),
    .A1(_04808_),
    .S(_04456_),
    .X(_05313_));
 sky130_fd_sc_hd__a21o_1 _11146_ (.A1(_01971_),
    .A2(_05313_),
    .B1(_04457_),
    .X(_05314_));
 sky130_fd_sc_hd__o221a_1 _11147_ (.A1(_02307_),
    .A2(_05308_),
    .B1(_05312_),
    .B2(_04790_),
    .C1(_05314_),
    .X(_05315_));
 sky130_fd_sc_hd__inv_2 _11148_ (.A(_04463_),
    .Y(_05316_));
 sky130_fd_sc_hd__o211a_1 _11149_ (.A1(_05316_),
    .A2(_05269_),
    .B1(_04458_),
    .C1(_04462_),
    .X(_05317_));
 sky130_fd_sc_hd__a21o_1 _11150_ (.A1(_01747_),
    .A2(_04466_),
    .B1(_04494_),
    .X(_05318_));
 sky130_fd_sc_hd__or2_1 _11151_ (.A(_04456_),
    .B(_04457_),
    .X(_05319_));
 sky130_fd_sc_hd__o211a_1 _11152_ (.A1(_05254_),
    .A2(_05318_),
    .B1(_05319_),
    .C1(_04463_),
    .X(_05320_));
 sky130_fd_sc_hd__a21oi_1 _11153_ (.A1(_05280_),
    .A2(_05266_),
    .B1(_05319_),
    .Y(_05321_));
 sky130_fd_sc_hd__a31o_1 _11154_ (.A1(_05319_),
    .A2(_05280_),
    .A3(_05266_),
    .B1(_04781_),
    .X(_05322_));
 sky130_fd_sc_hd__or2_1 _11155_ (.A(_05321_),
    .B(_05322_),
    .X(_05323_));
 sky130_fd_sc_hd__o311a_1 _11156_ (.A1(_04870_),
    .A2(_05317_),
    .A3(_05320_),
    .B1(_05323_),
    .C1(_04853_),
    .X(_05324_));
 sky130_fd_sc_hd__a21oi_1 _11157_ (.A1(_04402_),
    .A2(_05315_),
    .B1(_05324_),
    .Y(_05325_));
 sky130_fd_sc_hd__a211o_1 _11158_ (.A1(_05299_),
    .A2(_05300_),
    .B1(_05304_),
    .C1(_05325_),
    .X(_05326_));
 sky130_fd_sc_hd__a22o_1 _11159_ (.A1(_04742_),
    .A2(_05298_),
    .B1(_05326_),
    .B2(_04815_),
    .X(_05327_));
 sky130_fd_sc_hd__and2_2 _11160_ (.A(_04760_),
    .B(_05327_),
    .X(_05328_));
 sky130_fd_sc_hd__clkbuf_4 _11161_ (.A(_05328_),
    .X(_05329_));
 sky130_fd_sc_hd__mux2_1 _11162_ (.A0(_05329_),
    .A1(\regs[9][14] ),
    .S(_05188_),
    .X(_05330_));
 sky130_fd_sc_hd__clkbuf_1 _11163_ (.A(_05330_),
    .X(_00333_));
 sky130_fd_sc_hd__a221o_1 _11164_ (.A1(_02587_),
    .A2(_04183_),
    .B1(_05037_),
    .B2(_05036_),
    .C1(_05082_),
    .X(_05331_));
 sky130_fd_sc_hd__a21oi_2 _11165_ (.A1(_04945_),
    .A2(_05331_),
    .B1(_01984_),
    .Y(_05332_));
 sky130_fd_sc_hd__or3_1 _11166_ (.A(_04453_),
    .B(_04456_),
    .C(_05321_),
    .X(_05333_));
 sky130_fd_sc_hd__o21ai_1 _11167_ (.A1(_04456_),
    .A2(_05321_),
    .B1(_04453_),
    .Y(_05334_));
 sky130_fd_sc_hd__a21oi_1 _11168_ (.A1(_01871_),
    .A2(_04499_),
    .B1(_05320_),
    .Y(_05335_));
 sky130_fd_sc_hd__a21oi_1 _11169_ (.A1(_04453_),
    .A2(_05335_),
    .B1(_04870_),
    .Y(_05336_));
 sky130_fd_sc_hd__or2_1 _11170_ (.A(_04453_),
    .B(_05335_),
    .X(_05337_));
 sky130_fd_sc_hd__a32o_1 _11171_ (.A1(_04868_),
    .A2(_05333_),
    .A3(_05334_),
    .B1(_05336_),
    .B2(_05337_),
    .X(_05338_));
 sky130_fd_sc_hd__mux2_1 _11172_ (.A0(_05273_),
    .A1(_05281_),
    .S(_04622_),
    .X(_05339_));
 sky130_fd_sc_hd__o21a_1 _11173_ (.A1(_04926_),
    .A2(_05306_),
    .B1(_04879_),
    .X(_05340_));
 sky130_fd_sc_hd__o21ai_1 _11174_ (.A1(_04882_),
    .A2(_05339_),
    .B1(_05340_),
    .Y(_05341_));
 sky130_fd_sc_hd__o21a_1 _11175_ (.A1(_04926_),
    .A2(_05339_),
    .B1(_04879_),
    .X(_05342_));
 sky130_fd_sc_hd__o21ai_1 _11176_ (.A1(_04882_),
    .A2(_05310_),
    .B1(_05342_),
    .Y(_05343_));
 sky130_fd_sc_hd__or2_1 _11177_ (.A(_01870_),
    .B(_04452_),
    .X(_05344_));
 sky130_fd_sc_hd__a31o_1 _11178_ (.A1(_01870_),
    .A2(_04891_),
    .A3(_04452_),
    .B1(_04177_),
    .X(_05345_));
 sky130_fd_sc_hd__a221o_1 _11179_ (.A1(_05057_),
    .A2(_05344_),
    .B1(_04453_),
    .B2(_04831_),
    .C1(_05345_),
    .X(_05346_));
 sky130_fd_sc_hd__o21ba_1 _11180_ (.A1(_04933_),
    .A2(_05343_),
    .B1_N(_05346_),
    .X(_05347_));
 sky130_fd_sc_hd__o21ai_1 _11181_ (.A1(_02308_),
    .A2(_05341_),
    .B1(_05347_),
    .Y(_05348_));
 sky130_fd_sc_hd__o21ai_1 _11182_ (.A1(_04864_),
    .A2(_05338_),
    .B1(_05348_),
    .Y(_05349_));
 sky130_fd_sc_hd__or3_1 _11183_ (.A(_01613_),
    .B(_01618_),
    .C(_01622_),
    .X(_05350_));
 sky130_fd_sc_hd__o21ai_1 _11184_ (.A1(_01613_),
    .A2(_01622_),
    .B1(_01618_),
    .Y(_05351_));
 sky130_fd_sc_hd__buf_2 _11185_ (.A(_05227_),
    .X(_05352_));
 sky130_fd_sc_hd__a22o_1 _11186_ (.A1(\cycles[15] ),
    .A2(_05073_),
    .B1(_04390_),
    .B2(\cycles[47] ),
    .X(_05353_));
 sky130_fd_sc_hd__a221o_1 _11187_ (.A1(\instret[15] ),
    .A2(_04385_),
    .B1(_05072_),
    .B2(\instret[47] ),
    .C1(_05353_),
    .X(_05354_));
 sky130_fd_sc_hd__a22o_1 _11188_ (.A1(\J_type_imm[15] ),
    .A2(_05352_),
    .B1(_04376_),
    .B2(_05354_),
    .X(_05355_));
 sky130_fd_sc_hd__a31oi_1 _11189_ (.A1(_05299_),
    .A2(_05350_),
    .A3(_05351_),
    .B1(_05355_),
    .Y(_05356_));
 sky130_fd_sc_hd__o2111a_1 _11190_ (.A1(_01860_),
    .A2(_02071_),
    .B1(_05349_),
    .C1(_05356_),
    .D1(_01984_),
    .X(_05357_));
 sky130_fd_sc_hd__nor3_4 _11191_ (.A(_05032_),
    .B(_05332_),
    .C(_05357_),
    .Y(_05358_));
 sky130_fd_sc_hd__buf_2 _11192_ (.A(_05358_),
    .X(_05359_));
 sky130_fd_sc_hd__mux2_1 _11193_ (.A0(_05359_),
    .A1(\regs[9][15] ),
    .S(_05188_),
    .X(_05360_));
 sky130_fd_sc_hd__clkbuf_1 _11194_ (.A(_05360_),
    .X(_00334_));
 sky130_fd_sc_hd__nand2_1 _11195_ (.A(_04453_),
    .B(_04458_),
    .Y(_05361_));
 sky130_fd_sc_hd__a211o_1 _11196_ (.A1(_04462_),
    .A2(_04463_),
    .B1(_04468_),
    .C1(_05361_),
    .X(_05362_));
 sky130_fd_sc_hd__a21oi_1 _11197_ (.A1(_01872_),
    .A2(_04461_),
    .B1(_04465_),
    .Y(_05363_));
 sky130_fd_sc_hd__nand2_1 _11198_ (.A(_05344_),
    .B(_04456_),
    .Y(_05364_));
 sky130_fd_sc_hd__nand2_1 _11199_ (.A(_01870_),
    .B(_04452_),
    .Y(_05365_));
 sky130_fd_sc_hd__o311a_1 _11200_ (.A1(_05272_),
    .A2(_05361_),
    .A3(_05363_),
    .B1(_05364_),
    .C1(_05365_),
    .X(_05366_));
 sky130_fd_sc_hd__o21ai_1 _11201_ (.A1(_05249_),
    .A2(_05362_),
    .B1(_05366_),
    .Y(_05367_));
 sky130_fd_sc_hd__nor2_1 _11202_ (.A(_04525_),
    .B(_05367_),
    .Y(_05368_));
 sky130_fd_sc_hd__and2_1 _11203_ (.A(_04525_),
    .B(_05367_),
    .X(_05369_));
 sky130_fd_sc_hd__nor2_1 _11204_ (.A(_05368_),
    .B(_05369_),
    .Y(_05370_));
 sky130_fd_sc_hd__a311o_1 _11205_ (.A1(_04448_),
    .A2(_05067_),
    .A3(_05016_),
    .B1(_04404_),
    .C1(_04489_),
    .X(_05371_));
 sky130_fd_sc_hd__and3b_1 _11206_ (.A_N(_04459_),
    .B(_04463_),
    .C(_05318_),
    .X(_05372_));
 sky130_fd_sc_hd__a311oi_2 _11207_ (.A1(_01871_),
    .A2(_04500_),
    .A3(_04499_),
    .B1(_05372_),
    .C1(_04496_),
    .Y(_05373_));
 sky130_fd_sc_hd__nand2_1 _11208_ (.A(_04477_),
    .B(_05253_),
    .Y(_05374_));
 sky130_fd_sc_hd__o31a_1 _11209_ (.A1(_04479_),
    .A2(_04486_),
    .A3(_05175_),
    .B1(_05374_),
    .X(_05375_));
 sky130_fd_sc_hd__or2_1 _11210_ (.A(_04469_),
    .B(_05375_),
    .X(_05376_));
 sky130_fd_sc_hd__and3_1 _11211_ (.A(_05371_),
    .B(_05373_),
    .C(_05376_),
    .X(_05377_));
 sky130_fd_sc_hd__nand2_1 _11212_ (.A(_04525_),
    .B(_05377_),
    .Y(_05378_));
 sky130_fd_sc_hd__nor2_1 _11213_ (.A(_04525_),
    .B(_05377_),
    .Y(_05379_));
 sky130_fd_sc_hd__nor2_1 _11214_ (.A(_04786_),
    .B(_05379_),
    .Y(_05380_));
 sky130_fd_sc_hd__o211a_1 _11215_ (.A1(_04365_),
    .A2(_05370_),
    .B1(_05378_),
    .C1(_05380_),
    .X(_05381_));
 sky130_fd_sc_hd__a211o_1 _11216_ (.A1(_04780_),
    .A2(_05370_),
    .B1(_05381_),
    .C1(_04402_),
    .X(_05382_));
 sky130_fd_sc_hd__mux2_1 _11217_ (.A0(_04723_),
    .A1(_04827_),
    .S(_04522_),
    .X(_05383_));
 sky130_fd_sc_hd__a21o_1 _11218_ (.A1(_01972_),
    .A2(_05383_),
    .B1(_04524_),
    .X(_05384_));
 sky130_fd_sc_hd__o221a_1 _11219_ (.A1(_04933_),
    .A2(_05341_),
    .B1(_05343_),
    .B2(_04917_),
    .C1(_05384_),
    .X(_05385_));
 sky130_fd_sc_hd__nand2_1 _11220_ (.A(_04402_),
    .B(_05385_),
    .Y(_05386_));
 sky130_fd_sc_hd__xnor2_1 _11221_ (.A(_01557_),
    .B(_01623_),
    .Y(_05387_));
 sky130_fd_sc_hd__a22o_1 _11222_ (.A1(\cycles[16] ),
    .A2(_04391_),
    .B1(_04389_),
    .B2(\cycles[48] ),
    .X(_05388_));
 sky130_fd_sc_hd__a221o_2 _11223_ (.A1(\instret[16] ),
    .A2(_04384_),
    .B1(_04897_),
    .B2(\instret[48] ),
    .C1(_05388_),
    .X(_05389_));
 sky130_fd_sc_hd__a22o_1 _11224_ (.A1(\J_type_imm[16] ),
    .A2(_05227_),
    .B1(_04375_),
    .B2(_05389_),
    .X(_05390_));
 sky130_fd_sc_hd__nor2_1 _11225_ (.A(_01859_),
    .B(_02055_),
    .Y(_05391_));
 sky130_fd_sc_hd__a211o_1 _11226_ (.A1(_04863_),
    .A2(_05387_),
    .B1(_05390_),
    .C1(_05391_),
    .X(_05392_));
 sky130_fd_sc_hd__a311o_1 _11227_ (.A1(_04366_),
    .A2(_05382_),
    .A3(_05386_),
    .B1(_05392_),
    .C1(_01528_),
    .X(_05393_));
 sky130_fd_sc_hd__or2_1 _11228_ (.A(net8),
    .B(_04033_),
    .X(_05394_));
 sky130_fd_sc_hd__a41o_2 _11229_ (.A1(_01688_),
    .A2(_05036_),
    .A3(_05394_),
    .A4(_05034_),
    .B1(_05082_),
    .X(_05395_));
 sky130_fd_sc_hd__buf_2 _11230_ (.A(_05395_),
    .X(_05396_));
 sky130_fd_sc_hd__a21o_1 _11231_ (.A1(_02297_),
    .A2(_05033_),
    .B1(_05396_),
    .X(_05397_));
 sky130_fd_sc_hd__a21o_1 _11232_ (.A1(_04945_),
    .A2(_05397_),
    .B1(_04949_),
    .X(_05398_));
 sky130_fd_sc_hd__and3_2 _11233_ (.A(_04759_),
    .B(_05393_),
    .C(_05398_),
    .X(_05399_));
 sky130_fd_sc_hd__clkbuf_4 _11234_ (.A(_05399_),
    .X(_05400_));
 sky130_fd_sc_hd__mux2_1 _11235_ (.A0(_05400_),
    .A1(\regs[9][16] ),
    .S(_05188_),
    .X(_05401_));
 sky130_fd_sc_hd__clkbuf_1 _11236_ (.A(_05401_),
    .X(_00335_));
 sky130_fd_sc_hd__a21o_1 _11237_ (.A1(net10),
    .A2(_04733_),
    .B1(_05395_),
    .X(_05402_));
 sky130_fd_sc_hd__xnor2_1 _11238_ (.A(_01554_),
    .B(_01624_),
    .Y(_05403_));
 sky130_fd_sc_hd__a22o_1 _11239_ (.A1(\cycles[17] ),
    .A2(_04392_),
    .B1(_04389_),
    .B2(\cycles[49] ),
    .X(_05404_));
 sky130_fd_sc_hd__a221o_1 _11240_ (.A1(\instret[17] ),
    .A2(_04384_),
    .B1(_04395_),
    .B2(\instret[49] ),
    .C1(_05404_),
    .X(_05405_));
 sky130_fd_sc_hd__a22o_1 _11241_ (.A1(\J_type_imm[17] ),
    .A2(_05227_),
    .B1(_04375_),
    .B2(_05405_),
    .X(_05406_));
 sky130_fd_sc_hd__o21a_1 _11242_ (.A1(_04522_),
    .A2(_05369_),
    .B1(_04519_),
    .X(_05407_));
 sky130_fd_sc_hd__nor3_1 _11243_ (.A(_04519_),
    .B(_04522_),
    .C(_05369_),
    .Y(_05408_));
 sky130_fd_sc_hd__or3_1 _11244_ (.A(_04782_),
    .B(_05407_),
    .C(_05408_),
    .X(_05409_));
 sky130_fd_sc_hd__a21oi_1 _11245_ (.A1(_01868_),
    .A2(_04521_),
    .B1(_05379_),
    .Y(_05410_));
 sky130_fd_sc_hd__o21ai_1 _11246_ (.A1(_04519_),
    .A2(_05410_),
    .B1(_04787_),
    .Y(_05411_));
 sky130_fd_sc_hd__a21o_1 _11247_ (.A1(_04519_),
    .A2(_05410_),
    .B1(_05411_),
    .X(_05412_));
 sky130_fd_sc_hd__or2_1 _11248_ (.A(_04789_),
    .B(_05308_),
    .X(_05413_));
 sky130_fd_sc_hd__and2_1 _11249_ (.A(_01723_),
    .B(_04516_),
    .X(_05414_));
 sky130_fd_sc_hd__or2_1 _11250_ (.A(_01723_),
    .B(_04516_),
    .X(_05415_));
 sky130_fd_sc_hd__a221o_1 _11251_ (.A1(_01827_),
    .A2(_05414_),
    .B1(_05415_),
    .B2(_05057_),
    .C1(_04177_),
    .X(_05416_));
 sky130_fd_sc_hd__a21oi_1 _11252_ (.A1(_04831_),
    .A2(_04519_),
    .B1(_05416_),
    .Y(_05417_));
 sky130_fd_sc_hd__o211a_1 _11253_ (.A1(_02306_),
    .A2(_05312_),
    .B1(_05413_),
    .C1(_05417_),
    .X(_05418_));
 sky130_fd_sc_hd__a31o_1 _11254_ (.A1(_04853_),
    .A2(_05409_),
    .A3(_05412_),
    .B1(_05418_),
    .X(_05419_));
 sky130_fd_sc_hd__o21ai_1 _11255_ (.A1(_01859_),
    .A2(_02043_),
    .B1(_05419_),
    .Y(_05420_));
 sky130_fd_sc_hd__a211o_1 _11256_ (.A1(_05299_),
    .A2(_05403_),
    .B1(_05406_),
    .C1(_05420_),
    .X(_05421_));
 sky130_fd_sc_hd__a22o_1 _11257_ (.A1(_04742_),
    .A2(_05402_),
    .B1(_05421_),
    .B2(_04815_),
    .X(_05422_));
 sky130_fd_sc_hd__and2_2 _11258_ (.A(_04760_),
    .B(_05422_),
    .X(_05423_));
 sky130_fd_sc_hd__clkbuf_4 _11259_ (.A(_05423_),
    .X(_05424_));
 sky130_fd_sc_hd__mux2_1 _11260_ (.A0(_05424_),
    .A1(\regs[9][17] ),
    .S(_05188_),
    .X(_05425_));
 sky130_fd_sc_hd__clkbuf_1 _11261_ (.A(_05425_),
    .X(_00336_));
 sky130_fd_sc_hd__nor2_1 _11262_ (.A(_01860_),
    .B(_02029_),
    .Y(_05426_));
 sky130_fd_sc_hd__a22o_1 _11263_ (.A1(\cycles[18] ),
    .A2(_04392_),
    .B1(_04939_),
    .B2(\cycles[50] ),
    .X(_05427_));
 sky130_fd_sc_hd__a221o_1 _11264_ (.A1(\instret[18] ),
    .A2(_04896_),
    .B1(_04395_),
    .B2(\instret[50] ),
    .C1(_05427_),
    .X(_05428_));
 sky130_fd_sc_hd__a221o_1 _11265_ (.A1(\J_type_imm[18] ),
    .A2(_05352_),
    .B1(_04938_),
    .B2(_05428_),
    .C1(_01527_),
    .X(_05429_));
 sky130_fd_sc_hd__o21ba_1 _11266_ (.A1(_01552_),
    .A2(_01624_),
    .B1_N(_01553_),
    .X(_05430_));
 sky130_fd_sc_hd__o21ai_1 _11267_ (.A1(_01551_),
    .A2(_05430_),
    .B1(_04825_),
    .Y(_05431_));
 sky130_fd_sc_hd__a21oi_1 _11268_ (.A1(_01551_),
    .A2(_05430_),
    .B1(_05431_),
    .Y(_05432_));
 sky130_fd_sc_hd__o21ai_1 _11269_ (.A1(_01799_),
    .A2(_04523_),
    .B1(_04517_),
    .Y(_05433_));
 sky130_fd_sc_hd__o211a_1 _11270_ (.A1(_05379_),
    .A2(_05433_),
    .B1(_04507_),
    .C1(_04518_),
    .X(_05434_));
 sky130_fd_sc_hd__inv_2 _11271_ (.A(_04518_),
    .Y(_05435_));
 sky130_fd_sc_hd__nor2_1 _11272_ (.A(_04505_),
    .B(_04506_),
    .Y(_05436_));
 sky130_fd_sc_hd__o211a_1 _11273_ (.A1(_05435_),
    .A2(_05410_),
    .B1(_05436_),
    .C1(_04517_),
    .X(_05437_));
 sky130_fd_sc_hd__o31a_1 _11274_ (.A1(_04786_),
    .A2(_05434_),
    .A3(_05437_),
    .B1(_04866_),
    .X(_05438_));
 sky130_fd_sc_hd__o21a_1 _11275_ (.A1(_05414_),
    .A2(_05407_),
    .B1(_05436_),
    .X(_05439_));
 sky130_fd_sc_hd__or3_1 _11276_ (.A(_05436_),
    .B(_05414_),
    .C(_05407_),
    .X(_05440_));
 sky130_fd_sc_hd__or3b_1 _11277_ (.A(_05438_),
    .B(_05439_),
    .C_N(_05440_),
    .X(_05441_));
 sky130_fd_sc_hd__o31a_1 _11278_ (.A1(_04870_),
    .A2(_05434_),
    .A3(_05437_),
    .B1(_04178_),
    .X(_05442_));
 sky130_fd_sc_hd__nand2_1 _11279_ (.A(_01827_),
    .B(_04505_),
    .Y(_05443_));
 sky130_fd_sc_hd__o211a_1 _11280_ (.A1(_01829_),
    .A2(_04505_),
    .B1(_05443_),
    .C1(_01816_),
    .X(_05444_));
 sky130_fd_sc_hd__o22a_1 _11281_ (.A1(_02306_),
    .A2(_05276_),
    .B1(_05444_),
    .B2(_04506_),
    .X(_05445_));
 sky130_fd_sc_hd__o211a_1 _11282_ (.A1(_04790_),
    .A2(_05284_),
    .B1(_05445_),
    .C1(_04401_),
    .X(_05446_));
 sky130_fd_sc_hd__a211o_1 _11283_ (.A1(_05441_),
    .A2(_05442_),
    .B1(_05446_),
    .C1(_04728_),
    .X(_05447_));
 sky130_fd_sc_hd__or4b_1 _11284_ (.A(_05426_),
    .B(_05429_),
    .C(_05432_),
    .D_N(_05447_),
    .X(_05448_));
 sky130_fd_sc_hd__a21o_1 _11285_ (.A1(net11),
    .A2(_05033_),
    .B1(_05396_),
    .X(_05449_));
 sky130_fd_sc_hd__a21o_1 _11286_ (.A1(_04741_),
    .A2(_05449_),
    .B1(_04949_),
    .X(_05450_));
 sky130_fd_sc_hd__and3_2 _11287_ (.A(_04759_),
    .B(_05448_),
    .C(_05450_),
    .X(_05451_));
 sky130_fd_sc_hd__buf_2 _11288_ (.A(_05451_),
    .X(_05452_));
 sky130_fd_sc_hd__mux2_1 _11289_ (.A0(_05452_),
    .A1(\regs[9][18] ),
    .S(_05188_),
    .X(_05453_));
 sky130_fd_sc_hd__clkbuf_1 _11290_ (.A(_05453_),
    .X(_00337_));
 sky130_fd_sc_hd__a21o_1 _11291_ (.A1(net12),
    .A2(_04733_),
    .B1(_05395_),
    .X(_05454_));
 sky130_fd_sc_hd__a21o_1 _11292_ (.A1(_01550_),
    .A2(_05430_),
    .B1(_01549_),
    .X(_05455_));
 sky130_fd_sc_hd__xnor2_1 _11293_ (.A(_01630_),
    .B(_05455_),
    .Y(_05456_));
 sky130_fd_sc_hd__a22o_1 _11294_ (.A1(\cycles[19] ),
    .A2(_04392_),
    .B1(_04389_),
    .B2(\cycles[51] ),
    .X(_05457_));
 sky130_fd_sc_hd__a221o_1 _11295_ (.A1(\instret[19] ),
    .A2(_04384_),
    .B1(_04897_),
    .B2(\instret[51] ),
    .C1(_05457_),
    .X(_05458_));
 sky130_fd_sc_hd__a22oi_1 _11296_ (.A1(\J_type_imm[19] ),
    .A2(_05227_),
    .B1(_04375_),
    .B2(_05458_),
    .Y(_05459_));
 sky130_fd_sc_hd__o21ai_1 _11297_ (.A1(_01859_),
    .A2(_02018_),
    .B1(_05459_),
    .Y(_05460_));
 sky130_fd_sc_hd__or2_1 _11298_ (.A(_04511_),
    .B(_04512_),
    .X(_05461_));
 sky130_fd_sc_hd__o21ai_1 _11299_ (.A1(_04505_),
    .A2(_05439_),
    .B1(_05461_),
    .Y(_05462_));
 sky130_fd_sc_hd__or3_1 _11300_ (.A(_04505_),
    .B(_05461_),
    .C(_05439_),
    .X(_05463_));
 sky130_fd_sc_hd__o21ba_1 _11301_ (.A1(_04551_),
    .A2(_04504_),
    .B1_N(_05434_),
    .X(_05464_));
 sky130_fd_sc_hd__xnor2_1 _11302_ (.A(_04513_),
    .B(_05464_),
    .Y(_05465_));
 sky130_fd_sc_hd__a32o_1 _11303_ (.A1(_04867_),
    .A2(_05462_),
    .A3(_05463_),
    .B1(_05465_),
    .B2(_04787_),
    .X(_05466_));
 sky130_fd_sc_hd__nor2_1 _11304_ (.A(_04791_),
    .B(_05242_),
    .Y(_05467_));
 sky130_fd_sc_hd__nor2_1 _11305_ (.A(_02306_),
    .B(_05238_),
    .Y(_05468_));
 sky130_fd_sc_hd__or2_1 _11306_ (.A(_01717_),
    .B(_04509_),
    .X(_05469_));
 sky130_fd_sc_hd__and2_1 _11307_ (.A(_01717_),
    .B(_04509_),
    .X(_05470_));
 sky130_fd_sc_hd__a221o_1 _11308_ (.A1(_05057_),
    .A2(_05469_),
    .B1(_05470_),
    .B2(_04891_),
    .C1(_04177_),
    .X(_05471_));
 sky130_fd_sc_hd__a211o_1 _11309_ (.A1(_04831_),
    .A2(_05461_),
    .B1(_05468_),
    .C1(_05471_),
    .X(_05472_));
 sky130_fd_sc_hd__o22a_1 _11310_ (.A1(_04864_),
    .A2(_05466_),
    .B1(_05467_),
    .B2(_05472_),
    .X(_05473_));
 sky130_fd_sc_hd__a211o_1 _11311_ (.A1(_04863_),
    .A2(_05456_),
    .B1(_05460_),
    .C1(_05473_),
    .X(_05474_));
 sky130_fd_sc_hd__a22o_1 _11312_ (.A1(_04742_),
    .A2(_05454_),
    .B1(_05474_),
    .B2(_04815_),
    .X(_05475_));
 sky130_fd_sc_hd__and2_2 _11313_ (.A(_04760_),
    .B(_05475_),
    .X(_05476_));
 sky130_fd_sc_hd__buf_4 _11314_ (.A(_05476_),
    .X(_05477_));
 sky130_fd_sc_hd__mux2_1 _11315_ (.A0(_05477_),
    .A1(\regs[9][19] ),
    .S(_05188_),
    .X(_05478_));
 sky130_fd_sc_hd__clkbuf_1 _11316_ (.A(_05478_),
    .X(_00338_));
 sky130_fd_sc_hd__nor2_1 _11317_ (.A(_04917_),
    .B(_05201_),
    .Y(_05479_));
 sky130_fd_sc_hd__mux2_1 _11318_ (.A0(_04723_),
    .A1(_04827_),
    .S(_04543_),
    .X(_05480_));
 sky130_fd_sc_hd__a21oi_1 _11319_ (.A1(_01972_),
    .A2(_05480_),
    .B1(_04542_),
    .Y(_05481_));
 sky130_fd_sc_hd__nor2_1 _11320_ (.A(_04933_),
    .B(_05208_),
    .Y(_05482_));
 sky130_fd_sc_hd__o31a_1 _11321_ (.A1(_05479_),
    .A2(_05481_),
    .A3(_05482_),
    .B1(_04864_),
    .X(_05483_));
 sky130_fd_sc_hd__a22o_1 _11322_ (.A1(\cycles[20] ),
    .A2(_04391_),
    .B1(_04389_),
    .B2(\cycles[52] ),
    .X(_05484_));
 sky130_fd_sc_hd__a221o_1 _11323_ (.A1(\instret[20] ),
    .A2(_04384_),
    .B1(_04897_),
    .B2(\instret[52] ),
    .C1(_05484_),
    .X(_05485_));
 sky130_fd_sc_hd__xnor2_1 _11324_ (.A(_01546_),
    .B(\I_type_imm[0] ),
    .Y(_05486_));
 sky130_fd_sc_hd__a21boi_1 _11325_ (.A1(_01629_),
    .A2(_05455_),
    .B1_N(_01548_),
    .Y(_05487_));
 sky130_fd_sc_hd__nor2_1 _11326_ (.A(_05486_),
    .B(_05487_),
    .Y(_05488_));
 sky130_fd_sc_hd__nand2_1 _11327_ (.A(_05486_),
    .B(_05487_),
    .Y(_05489_));
 sky130_fd_sc_hd__and3b_1 _11328_ (.A_N(_05488_),
    .B(_04370_),
    .C(_05489_),
    .X(_05490_));
 sky130_fd_sc_hd__a221o_1 _11329_ (.A1(_01564_),
    .A2(_05227_),
    .B1(_04375_),
    .B2(_05485_),
    .C1(_05490_),
    .X(_05491_));
 sky130_fd_sc_hd__o21bai_1 _11330_ (.A1(_01860_),
    .A2(_01999_),
    .B1_N(_05491_),
    .Y(_05492_));
 sky130_fd_sc_hd__nor2_1 _11331_ (.A(_04507_),
    .B(_04513_),
    .Y(_05493_));
 sky130_fd_sc_hd__and3_1 _11332_ (.A(_04519_),
    .B(_04525_),
    .C(_05493_),
    .X(_05494_));
 sky130_fd_sc_hd__o21a_1 _11333_ (.A1(_05414_),
    .A2(_04522_),
    .B1(_05415_),
    .X(_05495_));
 sky130_fd_sc_hd__a221o_1 _11334_ (.A1(_04505_),
    .A2(_05469_),
    .B1(_05493_),
    .B2(_05495_),
    .C1(_05470_),
    .X(_05496_));
 sky130_fd_sc_hd__a21oi_1 _11335_ (.A1(_05367_),
    .A2(_05494_),
    .B1(_05496_),
    .Y(_05497_));
 sky130_fd_sc_hd__and2_1 _11336_ (.A(_04544_),
    .B(_05497_),
    .X(_05498_));
 sky130_fd_sc_hd__nor2_1 _11337_ (.A(_04544_),
    .B(_05497_),
    .Y(_05499_));
 sky130_fd_sc_hd__or4b_1 _11338_ (.A(_05436_),
    .B(_05461_),
    .C(_05435_),
    .D_N(_05433_),
    .X(_05500_));
 sky130_fd_sc_hd__o311a_1 _11339_ (.A1(_04551_),
    .A2(_04504_),
    .A3(_04512_),
    .B1(_05500_),
    .C1(_04510_),
    .X(_05501_));
 sky130_fd_sc_hd__o41a_1 _11340_ (.A1(_04514_),
    .A2(_04519_),
    .A3(_04525_),
    .A4(_05377_),
    .B1(_05501_),
    .X(_05502_));
 sky130_fd_sc_hd__and2_1 _11341_ (.A(_04545_),
    .B(_05502_),
    .X(_05503_));
 sky130_fd_sc_hd__nor2_1 _11342_ (.A(_04545_),
    .B(_05502_),
    .Y(_05504_));
 sky130_fd_sc_hd__nor2_1 _11343_ (.A(_05503_),
    .B(_05504_),
    .Y(_05505_));
 sky130_fd_sc_hd__a2bb2o_1 _11344_ (.A1_N(_05498_),
    .A2_N(_05499_),
    .B1(_05070_),
    .B2(_05505_),
    .X(_05506_));
 sky130_fd_sc_hd__inv_2 _11345_ (.A(_04786_),
    .Y(_05507_));
 sky130_fd_sc_hd__a21o_1 _11346_ (.A1(_05507_),
    .A2(_05505_),
    .B1(_04780_),
    .X(_05508_));
 sky130_fd_sc_hd__and4_1 _11347_ (.A(_04178_),
    .B(_04366_),
    .C(_05506_),
    .D(_05508_),
    .X(_05509_));
 sky130_fd_sc_hd__a21o_1 _11348_ (.A1(_03386_),
    .A2(_04182_),
    .B1(_05395_),
    .X(_05510_));
 sky130_fd_sc_hd__a21o_1 _11349_ (.A1(_04741_),
    .A2(_05510_),
    .B1(\core_state[1] ),
    .X(_05511_));
 sky130_fd_sc_hd__o41a_1 _11350_ (.A1(_01528_),
    .A2(_05483_),
    .A3(_05492_),
    .A4(_05509_),
    .B1(_05511_),
    .X(_05512_));
 sky130_fd_sc_hd__and2_2 _11351_ (.A(_04760_),
    .B(_05512_),
    .X(_05513_));
 sky130_fd_sc_hd__clkbuf_4 _11352_ (.A(_05513_),
    .X(_05514_));
 sky130_fd_sc_hd__buf_8 _11353_ (.A(_04768_),
    .X(_05515_));
 sky130_fd_sc_hd__mux2_1 _11354_ (.A0(_05514_),
    .A1(\regs[9][20] ),
    .S(_05515_),
    .X(_05516_));
 sky130_fd_sc_hd__clkbuf_1 _11355_ (.A(_05516_),
    .X(_00339_));
 sky130_fd_sc_hd__a21o_1 _11356_ (.A1(_02276_),
    .A2(_04733_),
    .B1(_05395_),
    .X(_05517_));
 sky130_fd_sc_hd__or2_1 _11357_ (.A(\PC[21] ),
    .B(_02275_),
    .X(_05518_));
 sky130_fd_sc_hd__nand2_1 _11358_ (.A(\PC[21] ),
    .B(_02275_),
    .Y(_05519_));
 sky130_fd_sc_hd__nand2_1 _11359_ (.A(_05518_),
    .B(_05519_),
    .Y(_05520_));
 sky130_fd_sc_hd__a21o_1 _11360_ (.A1(_01546_),
    .A2(_01564_),
    .B1(_05488_),
    .X(_05521_));
 sky130_fd_sc_hd__xnor2_1 _11361_ (.A(_05520_),
    .B(_05521_),
    .Y(_05522_));
 sky130_fd_sc_hd__nor2_1 _11362_ (.A(_01859_),
    .B(_01995_),
    .Y(_05523_));
 sky130_fd_sc_hd__a22o_1 _11363_ (.A1(\cycles[21] ),
    .A2(_04392_),
    .B1(_04389_),
    .B2(\cycles[53] ),
    .X(_05524_));
 sky130_fd_sc_hd__a221o_1 _11364_ (.A1(\instret[21] ),
    .A2(_04384_),
    .B1(_04897_),
    .B2(\instret[53] ),
    .C1(_05524_),
    .X(_05525_));
 sky130_fd_sc_hd__a22o_1 _11365_ (.A1(_02275_),
    .A2(_05227_),
    .B1(_04375_),
    .B2(_05525_),
    .X(_05526_));
 sky130_fd_sc_hd__o21ai_1 _11366_ (.A1(_04543_),
    .A2(_05499_),
    .B1(_04540_),
    .Y(_05527_));
 sky130_fd_sc_hd__o311a_1 _11367_ (.A1(_04540_),
    .A2(_04543_),
    .A3(_05499_),
    .B1(_05527_),
    .C1(_04867_),
    .X(_05528_));
 sky130_fd_sc_hd__a21o_1 _11368_ (.A1(\leorv32_alu.input1[20] ),
    .A2(_04541_),
    .B1(_05504_),
    .X(_05529_));
 sky130_fd_sc_hd__or2_1 _11369_ (.A(_04540_),
    .B(_05529_),
    .X(_05530_));
 sky130_fd_sc_hd__nand2_1 _11370_ (.A(_04540_),
    .B(_05529_),
    .Y(_05531_));
 sky130_fd_sc_hd__a21oi_1 _11371_ (.A1(_05530_),
    .A2(_05531_),
    .B1(_04870_),
    .Y(_05532_));
 sky130_fd_sc_hd__nor2_1 _11372_ (.A(_04791_),
    .B(_05163_),
    .Y(_05533_));
 sky130_fd_sc_hd__nor2_1 _11373_ (.A(_02306_),
    .B(_05169_),
    .Y(_05534_));
 sky130_fd_sc_hd__a221o_1 _11374_ (.A1(_04891_),
    .A2(_04537_),
    .B1(_04539_),
    .B2(_05057_),
    .C1(_04177_),
    .X(_05535_));
 sky130_fd_sc_hd__a211o_1 _11375_ (.A1(_04831_),
    .A2(_04540_),
    .B1(_05534_),
    .C1(_05535_),
    .X(_05536_));
 sky130_fd_sc_hd__o32a_1 _11376_ (.A1(_04729_),
    .A2(_05528_),
    .A3(_05532_),
    .B1(_05533_),
    .B2(_05536_),
    .X(_05537_));
 sky130_fd_sc_hd__a2111o_1 _11377_ (.A1(_04863_),
    .A2(_05522_),
    .B1(_05523_),
    .C1(_05526_),
    .D1(_05537_),
    .X(_05538_));
 sky130_fd_sc_hd__a22o_1 _11378_ (.A1(_04742_),
    .A2(_05517_),
    .B1(_05538_),
    .B2(\core_state[1] ),
    .X(_05539_));
 sky130_fd_sc_hd__and2_1 _11379_ (.A(_04760_),
    .B(_05539_),
    .X(_05540_));
 sky130_fd_sc_hd__clkbuf_4 _11380_ (.A(_05540_),
    .X(_05541_));
 sky130_fd_sc_hd__mux2_1 _11381_ (.A0(_05541_),
    .A1(\regs[9][21] ),
    .S(_05515_),
    .X(_05542_));
 sky130_fd_sc_hd__clkbuf_1 _11382_ (.A(_05542_),
    .X(_00340_));
 sky130_fd_sc_hd__and2_1 _11383_ (.A(\PC[22] ),
    .B(_01900_),
    .X(_05543_));
 sky130_fd_sc_hd__nor2_1 _11384_ (.A(\PC[22] ),
    .B(_01900_),
    .Y(_05544_));
 sky130_fd_sc_hd__nor2_1 _11385_ (.A(_05543_),
    .B(_05544_),
    .Y(_05545_));
 sky130_fd_sc_hd__a221o_1 _11386_ (.A1(\PC[21] ),
    .A2(_02275_),
    .B1(_01564_),
    .B2(_01546_),
    .C1(_05488_),
    .X(_05546_));
 sky130_fd_sc_hd__and3_1 _11387_ (.A(_05518_),
    .B(_05545_),
    .C(_05546_),
    .X(_05547_));
 sky130_fd_sc_hd__and2_1 _11388_ (.A(_05518_),
    .B(_05546_),
    .X(_05548_));
 sky130_fd_sc_hd__o21ai_1 _11389_ (.A1(_05545_),
    .A2(_05548_),
    .B1(_05299_),
    .Y(_05549_));
 sky130_fd_sc_hd__a22o_1 _11390_ (.A1(\cycles[22] ),
    .A2(_04392_),
    .B1(_04939_),
    .B2(\cycles[54] ),
    .X(_05550_));
 sky130_fd_sc_hd__a221o_1 _11391_ (.A1(\instret[22] ),
    .A2(_04896_),
    .B1(_04395_),
    .B2(\instret[54] ),
    .C1(_05550_),
    .X(_05551_));
 sky130_fd_sc_hd__a22o_1 _11392_ (.A1(_01900_),
    .A2(_05352_),
    .B1(_04938_),
    .B2(_05551_),
    .X(_05552_));
 sky130_fd_sc_hd__o21ba_1 _11393_ (.A1(_01860_),
    .A2(_01974_),
    .B1_N(_05552_),
    .X(_05553_));
 sky130_fd_sc_hd__mux2_1 _11394_ (.A0(_04723_),
    .A1(_04827_),
    .S(_04527_),
    .X(_05554_));
 sky130_fd_sc_hd__a21o_1 _11395_ (.A1(_01972_),
    .A2(_05554_),
    .B1(_04529_),
    .X(_05555_));
 sky130_fd_sc_hd__o221a_1 _11396_ (.A1(_04917_),
    .A2(_05137_),
    .B1(_05143_),
    .B2(_04933_),
    .C1(_05555_),
    .X(_05556_));
 sky130_fd_sc_hd__or2_1 _11397_ (.A(_04527_),
    .B(_04529_),
    .X(_05557_));
 sky130_fd_sc_hd__a21oi_1 _11398_ (.A1(_04538_),
    .A2(_05527_),
    .B1(_05557_),
    .Y(_05558_));
 sky130_fd_sc_hd__a31o_1 _11399_ (.A1(_05557_),
    .A2(_04538_),
    .A3(_05527_),
    .B1(_04782_),
    .X(_05559_));
 sky130_fd_sc_hd__a211o_1 _11400_ (.A1(_04555_),
    .A2(_05529_),
    .B1(_04554_),
    .C1(_05557_),
    .X(_05560_));
 sky130_fd_sc_hd__a21o_1 _11401_ (.A1(\leorv32_alu.input1[20] ),
    .A2(_04541_),
    .B1(_04554_),
    .X(_05561_));
 sky130_fd_sc_hd__o211ai_2 _11402_ (.A1(_05561_),
    .A2(_05504_),
    .B1(_05557_),
    .C1(_04555_),
    .Y(_05562_));
 sky130_fd_sc_hd__a31o_1 _11403_ (.A1(_05070_),
    .A2(_05560_),
    .A3(_05562_),
    .B1(_04729_),
    .X(_05563_));
 sky130_fd_sc_hd__o21ba_1 _11404_ (.A1(_05558_),
    .A2(_05559_),
    .B1_N(_05563_),
    .X(_05564_));
 sky130_fd_sc_hd__a21o_1 _11405_ (.A1(_04402_),
    .A2(_05556_),
    .B1(_05564_),
    .X(_05565_));
 sky130_fd_sc_hd__o211ai_1 _11406_ (.A1(_05547_),
    .A2(_05549_),
    .B1(_05553_),
    .C1(_05565_),
    .Y(_05566_));
 sky130_fd_sc_hd__a21o_1 _11407_ (.A1(net16),
    .A2(_04183_),
    .B1(_05396_),
    .X(_05567_));
 sky130_fd_sc_hd__a21o_1 _11408_ (.A1(_04945_),
    .A2(_05567_),
    .B1(_01984_),
    .X(_05568_));
 sky130_fd_sc_hd__o211a_1 _11409_ (.A1(_01528_),
    .A2(_05566_),
    .B1(_05568_),
    .C1(_04771_),
    .X(_05569_));
 sky130_fd_sc_hd__clkbuf_4 _11410_ (.A(_05569_),
    .X(_05570_));
 sky130_fd_sc_hd__mux2_1 _11411_ (.A0(_05570_),
    .A1(\regs[9][22] ),
    .S(_05515_),
    .X(_05571_));
 sky130_fd_sc_hd__clkbuf_1 _11412_ (.A(_05571_),
    .X(_00341_));
 sky130_fd_sc_hd__nor2_1 _11413_ (.A(\PC[23] ),
    .B(_01897_),
    .Y(_05572_));
 sky130_fd_sc_hd__and2_1 _11414_ (.A(\PC[23] ),
    .B(_01897_),
    .X(_05573_));
 sky130_fd_sc_hd__nor2_1 _11415_ (.A(_05572_),
    .B(_05573_),
    .Y(_05574_));
 sky130_fd_sc_hd__or2_1 _11416_ (.A(_05543_),
    .B(_05547_),
    .X(_05575_));
 sky130_fd_sc_hd__nand2_1 _11417_ (.A(_05574_),
    .B(_05575_),
    .Y(_05576_));
 sky130_fd_sc_hd__o21a_1 _11418_ (.A1(_05574_),
    .A2(_05575_),
    .B1(_05299_),
    .X(_05577_));
 sky130_fd_sc_hd__nor2_1 _11419_ (.A(_02308_),
    .B(_05098_),
    .Y(_05578_));
 sky130_fd_sc_hd__nor2_1 _11420_ (.A(_04791_),
    .B(_05090_),
    .Y(_05579_));
 sky130_fd_sc_hd__or2_1 _11421_ (.A(\leorv32_alu.input1[23] ),
    .B(_04531_),
    .X(_05580_));
 sky130_fd_sc_hd__and2_1 _11422_ (.A(\leorv32_alu.input1[23] ),
    .B(_04531_),
    .X(_05581_));
 sky130_fd_sc_hd__a221o_1 _11423_ (.A1(_05057_),
    .A2(_05580_),
    .B1(_05581_),
    .B2(_04891_),
    .C1(_04178_),
    .X(_05582_));
 sky130_fd_sc_hd__a211o_1 _11424_ (.A1(_04831_),
    .A2(_04534_),
    .B1(_05579_),
    .C1(_05582_),
    .X(_05583_));
 sky130_fd_sc_hd__or3_1 _11425_ (.A(_04527_),
    .B(_04534_),
    .C(_05558_),
    .X(_05584_));
 sky130_fd_sc_hd__o21ai_1 _11426_ (.A1(_04527_),
    .A2(_05558_),
    .B1(_04534_),
    .Y(_05585_));
 sky130_fd_sc_hd__nand2_1 _11427_ (.A(\leorv32_alu.input1[22] ),
    .B(_04526_),
    .Y(_05586_));
 sky130_fd_sc_hd__a21oi_1 _11428_ (.A1(_05586_),
    .A2(_05562_),
    .B1(_04534_),
    .Y(_05587_));
 sky130_fd_sc_hd__a31o_1 _11429_ (.A1(_05586_),
    .A2(_04534_),
    .A3(_05562_),
    .B1(_04850_),
    .X(_05588_));
 sky130_fd_sc_hd__o21ai_1 _11430_ (.A1(_05587_),
    .A2(_05588_),
    .B1(_04853_),
    .Y(_05589_));
 sky130_fd_sc_hd__a31o_1 _11431_ (.A1(_04868_),
    .A2(_05584_),
    .A3(_05585_),
    .B1(_05589_),
    .X(_05590_));
 sky130_fd_sc_hd__o21a_1 _11432_ (.A1(_05578_),
    .A2(_05583_),
    .B1(_05590_),
    .X(_05591_));
 sky130_fd_sc_hd__a22o_1 _11433_ (.A1(\cycles[23] ),
    .A2(_04393_),
    .B1(_04390_),
    .B2(\cycles[55] ),
    .X(_05592_));
 sky130_fd_sc_hd__a221o_1 _11434_ (.A1(\instret[23] ),
    .A2(_04385_),
    .B1(_05072_),
    .B2(\instret[55] ),
    .C1(_05592_),
    .X(_05593_));
 sky130_fd_sc_hd__a2bb2o_1 _11435_ (.A1_N(_01859_),
    .A2_N(_01852_),
    .B1(_05227_),
    .B2(_01897_),
    .X(_05594_));
 sky130_fd_sc_hd__a21o_1 _11436_ (.A1(_04376_),
    .A2(_05593_),
    .B1(_05594_),
    .X(_05595_));
 sky130_fd_sc_hd__a211o_1 _11437_ (.A1(_05576_),
    .A2(_05577_),
    .B1(_05591_),
    .C1(_05595_),
    .X(_05596_));
 sky130_fd_sc_hd__a21o_1 _11438_ (.A1(net17),
    .A2(_04183_),
    .B1(_05396_),
    .X(_05597_));
 sky130_fd_sc_hd__a21o_1 _11439_ (.A1(_04945_),
    .A2(_05597_),
    .B1(_04949_),
    .X(_05598_));
 sky130_fd_sc_hd__o211a_1 _11440_ (.A1(_01528_),
    .A2(_05596_),
    .B1(_05598_),
    .C1(_04771_),
    .X(_05599_));
 sky130_fd_sc_hd__buf_2 _11441_ (.A(_05599_),
    .X(_05600_));
 sky130_fd_sc_hd__mux2_1 _11442_ (.A0(_05600_),
    .A1(\regs[9][23] ),
    .S(_05515_),
    .X(_05601_));
 sky130_fd_sc_hd__clkbuf_1 _11443_ (.A(_05601_),
    .X(_00342_));
 sky130_fd_sc_hd__o2111ai_1 _11444_ (.A1(_04537_),
    .A2(_04543_),
    .B1(_04539_),
    .C1(_04530_),
    .D1(_04534_),
    .Y(_05602_));
 sky130_fd_sc_hd__inv_2 _11445_ (.A(_04540_),
    .Y(_05603_));
 sky130_fd_sc_hd__nand2_1 _11446_ (.A(_04530_),
    .B(_04534_),
    .Y(_05604_));
 sky130_fd_sc_hd__a21oi_1 _11447_ (.A1(_04527_),
    .A2(_05580_),
    .B1(_05581_),
    .Y(_05605_));
 sky130_fd_sc_hd__o41a_1 _11448_ (.A1(_05603_),
    .A2(_04544_),
    .A3(_05497_),
    .A4(_05604_),
    .B1(_05605_),
    .X(_05606_));
 sky130_fd_sc_hd__and2_1 _11449_ (.A(_05602_),
    .B(_05606_),
    .X(_05607_));
 sky130_fd_sc_hd__xor2_1 _11450_ (.A(_04567_),
    .B(_05607_),
    .X(_05608_));
 sky130_fd_sc_hd__or2_1 _11451_ (.A(_04546_),
    .B(_05501_),
    .X(_05609_));
 sky130_fd_sc_hd__a31o_1 _11452_ (.A1(_05371_),
    .A2(_05373_),
    .A3(_05376_),
    .B1(_04547_),
    .X(_05610_));
 sky130_fd_sc_hd__nand2_1 _11453_ (.A(_04555_),
    .B(_05561_),
    .Y(_05611_));
 sky130_fd_sc_hd__o221a_1 _11454_ (.A1(_05586_),
    .A2(_04557_),
    .B1(_04535_),
    .B2(_05611_),
    .C1(_04532_),
    .X(_05612_));
 sky130_fd_sc_hd__and3_1 _11455_ (.A(_05609_),
    .B(_05610_),
    .C(_05612_),
    .X(_05613_));
 sky130_fd_sc_hd__and2_1 _11456_ (.A(_04567_),
    .B(_05613_),
    .X(_05614_));
 sky130_fd_sc_hd__nor2_1 _11457_ (.A(_04567_),
    .B(_05613_),
    .Y(_05615_));
 sky130_fd_sc_hd__nor2_1 _11458_ (.A(_05614_),
    .B(_05615_),
    .Y(_05616_));
 sky130_fd_sc_hd__nand2_1 _11459_ (.A(_05070_),
    .B(_05616_),
    .Y(_05617_));
 sky130_fd_sc_hd__a21oi_1 _11460_ (.A1(_05507_),
    .A2(_05616_),
    .B1(_04780_),
    .Y(_05618_));
 sky130_fd_sc_hd__a21oi_2 _11461_ (.A1(_05608_),
    .A2(_05617_),
    .B1(_05618_),
    .Y(_05619_));
 sky130_fd_sc_hd__or2_1 _11462_ (.A(\PC[23] ),
    .B(_01897_),
    .X(_05620_));
 sky130_fd_sc_hd__o311a_1 _11463_ (.A1(_05543_),
    .A2(_05547_),
    .A3(_05573_),
    .B1(_05620_),
    .C1(_01892_),
    .X(_05621_));
 sky130_fd_sc_hd__o21a_1 _11464_ (.A1(_05573_),
    .A2(_05575_),
    .B1(_05620_),
    .X(_05622_));
 sky130_fd_sc_hd__o21ai_1 _11465_ (.A1(_01892_),
    .A2(_05622_),
    .B1(_04863_),
    .Y(_05623_));
 sky130_fd_sc_hd__mux2_1 _11466_ (.A0(_01829_),
    .A1(_04808_),
    .S(_04566_),
    .X(_05624_));
 sky130_fd_sc_hd__a21o_1 _11467_ (.A1(_01971_),
    .A2(_05624_),
    .B1(_04565_),
    .X(_05625_));
 sky130_fd_sc_hd__o221a_1 _11468_ (.A1(_04791_),
    .A2(_05048_),
    .B1(_05055_),
    .B2(_02307_),
    .C1(_05625_),
    .X(_05626_));
 sky130_fd_sc_hd__a22o_1 _11469_ (.A1(\cycles[24] ),
    .A2(_04391_),
    .B1(_04388_),
    .B2(\cycles[56] ),
    .X(_05627_));
 sky130_fd_sc_hd__a221o_1 _11470_ (.A1(\instret[24] ),
    .A2(_04383_),
    .B1(_04897_),
    .B2(\instret[56] ),
    .C1(_05627_),
    .X(_05628_));
 sky130_fd_sc_hd__a221o_1 _11471_ (.A1(_01892_),
    .A2(_05227_),
    .B1(_04374_),
    .B2(_05628_),
    .C1(_01526_),
    .X(_05629_));
 sky130_fd_sc_hd__o21ba_1 _11472_ (.A1(_04853_),
    .A2(_05626_),
    .B1_N(_05629_),
    .X(_05630_));
 sky130_fd_sc_hd__o21ai_1 _11473_ (.A1(_05621_),
    .A2(_05623_),
    .B1(_05630_),
    .Y(_05631_));
 sky130_fd_sc_hd__a31o_1 _11474_ (.A1(_04178_),
    .A2(_04366_),
    .A3(_05619_),
    .B1(_05631_),
    .X(_05632_));
 sky130_fd_sc_hd__a21o_1 _11475_ (.A1(net18),
    .A2(_05033_),
    .B1(_05396_),
    .X(_05633_));
 sky130_fd_sc_hd__a21o_1 _11476_ (.A1(_04741_),
    .A2(_05633_),
    .B1(_04949_),
    .X(_05634_));
 sky130_fd_sc_hd__and3_1 _11477_ (.A(_04759_),
    .B(_05632_),
    .C(_05634_),
    .X(_05635_));
 sky130_fd_sc_hd__buf_2 _11478_ (.A(_05635_),
    .X(_05636_));
 sky130_fd_sc_hd__mux2_1 _11479_ (.A0(_05636_),
    .A1(\regs[9][24] ),
    .S(_05515_),
    .X(_05637_));
 sky130_fd_sc_hd__clkbuf_1 _11480_ (.A(_05637_),
    .X(_00343_));
 sky130_fd_sc_hd__nand2_1 _11481_ (.A(_01890_),
    .B(_05621_),
    .Y(_05638_));
 sky130_fd_sc_hd__or2_1 _11482_ (.A(_01890_),
    .B(_05621_),
    .X(_05639_));
 sky130_fd_sc_hd__a22o_1 _11483_ (.A1(\cycles[25] ),
    .A2(_05073_),
    .B1(_04939_),
    .B2(\cycles[57] ),
    .X(_05640_));
 sky130_fd_sc_hd__a221o_1 _11484_ (.A1(\instret[25] ),
    .A2(_04896_),
    .B1(_04395_),
    .B2(\instret[57] ),
    .C1(_05640_),
    .X(_05641_));
 sky130_fd_sc_hd__a221o_1 _11485_ (.A1(_01890_),
    .A2(_05352_),
    .B1(_04938_),
    .B2(_05641_),
    .C1(_01527_),
    .X(_05642_));
 sky130_fd_sc_hd__a21boi_1 _11486_ (.A1(_05602_),
    .A2(_05606_),
    .B1_N(_04567_),
    .Y(_05643_));
 sky130_fd_sc_hd__or3_1 _11487_ (.A(_04563_),
    .B(_04566_),
    .C(_05643_),
    .X(_05644_));
 sky130_fd_sc_hd__o21a_1 _11488_ (.A1(_04566_),
    .A2(_05643_),
    .B1(_04563_),
    .X(_05645_));
 sky130_fd_sc_hd__nor2_1 _11489_ (.A(_04782_),
    .B(_05645_),
    .Y(_05646_));
 sky130_fd_sc_hd__nor2_1 _11490_ (.A(_01703_),
    .B(_04564_),
    .Y(_05647_));
 sky130_fd_sc_hd__or2_1 _11491_ (.A(_05647_),
    .B(_05615_),
    .X(_05648_));
 sky130_fd_sc_hd__xnor2_1 _11492_ (.A(_04563_),
    .B(_05648_),
    .Y(_05649_));
 sky130_fd_sc_hd__a22o_1 _11493_ (.A1(_05644_),
    .A2(_05646_),
    .B1(_05649_),
    .B2(_05070_),
    .X(_05650_));
 sky130_fd_sc_hd__nor2_1 _11494_ (.A(_02308_),
    .B(_05010_),
    .Y(_05651_));
 sky130_fd_sc_hd__nor2_1 _11495_ (.A(_04791_),
    .B(_05002_),
    .Y(_05652_));
 sky130_fd_sc_hd__a221o_1 _11496_ (.A1(_04891_),
    .A2(_04561_),
    .B1(_04562_),
    .B2(_05057_),
    .C1(_04178_),
    .X(_05653_));
 sky130_fd_sc_hd__a211o_1 _11497_ (.A1(_04831_),
    .A2(_04563_),
    .B1(_05652_),
    .C1(_05653_),
    .X(_05654_));
 sky130_fd_sc_hd__o22a_1 _11498_ (.A1(_04864_),
    .A2(_05650_),
    .B1(_05651_),
    .B2(_05654_),
    .X(_05655_));
 sky130_fd_sc_hd__a311o_1 _11499_ (.A1(_05299_),
    .A2(_05638_),
    .A3(_05639_),
    .B1(_05642_),
    .C1(_05655_),
    .X(_05656_));
 sky130_fd_sc_hd__a21o_1 _11500_ (.A1(net19),
    .A2(_05033_),
    .B1(_05396_),
    .X(_05657_));
 sky130_fd_sc_hd__a21o_1 _11501_ (.A1(_04741_),
    .A2(_05657_),
    .B1(_04949_),
    .X(_05658_));
 sky130_fd_sc_hd__and3_1 _11502_ (.A(_04759_),
    .B(_05656_),
    .C(_05658_),
    .X(_05659_));
 sky130_fd_sc_hd__buf_2 _11503_ (.A(_05659_),
    .X(_05660_));
 sky130_fd_sc_hd__mux2_1 _11504_ (.A0(_05660_),
    .A1(\regs[9][25] ),
    .S(_05515_),
    .X(_05661_));
 sky130_fd_sc_hd__clkbuf_1 _11505_ (.A(_05661_),
    .X(_00344_));
 sky130_fd_sc_hd__nor2_1 _11506_ (.A(_04561_),
    .B(_05645_),
    .Y(_05662_));
 sky130_fd_sc_hd__xnor2_1 _11507_ (.A(_04571_),
    .B(_05662_),
    .Y(_05663_));
 sky130_fd_sc_hd__or2_1 _11508_ (.A(_04601_),
    .B(_05647_),
    .X(_05664_));
 sky130_fd_sc_hd__o211a_1 _11509_ (.A1(_05615_),
    .A2(_05664_),
    .B1(_04571_),
    .C1(_04599_),
    .X(_05665_));
 sky130_fd_sc_hd__a211oi_1 _11510_ (.A1(_04599_),
    .A2(_05648_),
    .B1(_04601_),
    .C1(_04571_),
    .Y(_05666_));
 sky130_fd_sc_hd__o31a_1 _11511_ (.A1(_04870_),
    .A2(_05665_),
    .A3(_05666_),
    .B1(_04853_),
    .X(_05667_));
 sky130_fd_sc_hd__o21ai_2 _11512_ (.A1(_04782_),
    .A2(_05663_),
    .B1(_05667_),
    .Y(_05668_));
 sky130_fd_sc_hd__nor2_1 _11513_ (.A(_04917_),
    .B(_04978_),
    .Y(_05669_));
 sky130_fd_sc_hd__nor2_1 _11514_ (.A(_04933_),
    .B(_04970_),
    .Y(_05670_));
 sky130_fd_sc_hd__mux2_1 _11515_ (.A0(_04723_),
    .A1(_04827_),
    .S(_04569_),
    .X(_05671_));
 sky130_fd_sc_hd__a21oi_1 _11516_ (.A1(_01972_),
    .A2(_05671_),
    .B1(_04570_),
    .Y(_05672_));
 sky130_fd_sc_hd__or4_2 _11517_ (.A(_04178_),
    .B(_05669_),
    .C(_05670_),
    .D(_05672_),
    .X(_05673_));
 sky130_fd_sc_hd__a22o_1 _11518_ (.A1(\cycles[26] ),
    .A2(_05073_),
    .B1(_04939_),
    .B2(\cycles[58] ),
    .X(_05674_));
 sky130_fd_sc_hd__a221o_1 _11519_ (.A1(\instret[26] ),
    .A2(_04896_),
    .B1(_05072_),
    .B2(\instret[58] ),
    .C1(_05674_),
    .X(_05675_));
 sky130_fd_sc_hd__and3_1 _11520_ (.A(_01595_),
    .B(_01890_),
    .C(_05621_),
    .X(_05676_));
 sky130_fd_sc_hd__a21o_1 _11521_ (.A1(_01890_),
    .A2(_05621_),
    .B1(_01595_),
    .X(_05677_));
 sky130_fd_sc_hd__and3b_1 _11522_ (.A_N(_05676_),
    .B(_05677_),
    .C(_04825_),
    .X(_05678_));
 sky130_fd_sc_hd__a221o_1 _11523_ (.A1(_01595_),
    .A2(_05352_),
    .B1(_04938_),
    .B2(_05675_),
    .C1(_05678_),
    .X(_05679_));
 sky130_fd_sc_hd__a211o_1 _11524_ (.A1(_05668_),
    .A2(_05673_),
    .B1(_05679_),
    .C1(_01528_),
    .X(_05680_));
 sky130_fd_sc_hd__a21o_1 _11525_ (.A1(net20),
    .A2(_05033_),
    .B1(_05396_),
    .X(_05681_));
 sky130_fd_sc_hd__a21o_1 _11526_ (.A1(_04741_),
    .A2(_05681_),
    .B1(_04949_),
    .X(_05682_));
 sky130_fd_sc_hd__and3_1 _11527_ (.A(_04759_),
    .B(_05680_),
    .C(_05682_),
    .X(_05683_));
 sky130_fd_sc_hd__clkbuf_4 _11528_ (.A(_05683_),
    .X(_05684_));
 sky130_fd_sc_hd__mux2_1 _11529_ (.A0(_05684_),
    .A1(\regs[9][26] ),
    .S(_05515_),
    .X(_05685_));
 sky130_fd_sc_hd__clkbuf_1 _11530_ (.A(_05685_),
    .X(_00345_));
 sky130_fd_sc_hd__nor3_1 _11531_ (.A(_04569_),
    .B(_04561_),
    .C(_05645_),
    .Y(_05686_));
 sky130_fd_sc_hd__o21ai_1 _11532_ (.A1(_04570_),
    .A2(_05686_),
    .B1(_04576_),
    .Y(_05687_));
 sky130_fd_sc_hd__o31a_1 _11533_ (.A1(_04570_),
    .A2(_04576_),
    .A3(_05686_),
    .B1(_04868_),
    .X(_05688_));
 sky130_fd_sc_hd__a21o_1 _11534_ (.A1(\leorv32_alu.input1[26] ),
    .A2(_04568_),
    .B1(_05665_),
    .X(_05689_));
 sky130_fd_sc_hd__xnor2_1 _11535_ (.A(_04576_),
    .B(_05689_),
    .Y(_05690_));
 sky130_fd_sc_hd__o2bb2a_1 _11536_ (.A1_N(_05687_),
    .A2_N(_05688_),
    .B1(_05690_),
    .B2(_04870_),
    .X(_05691_));
 sky130_fd_sc_hd__nor2_1 _11537_ (.A(_01700_),
    .B(_04572_),
    .Y(_05692_));
 sky130_fd_sc_hd__nand2_1 _11538_ (.A(_01700_),
    .B(_04572_),
    .Y(_05693_));
 sky130_fd_sc_hd__a221o_1 _11539_ (.A1(_04891_),
    .A2(_05692_),
    .B1(_05693_),
    .B2(_05057_),
    .C1(_04178_),
    .X(_05694_));
 sky130_fd_sc_hd__o21ba_1 _11540_ (.A1(_01823_),
    .A2(_04576_),
    .B1_N(_05694_),
    .X(_05695_));
 sky130_fd_sc_hd__o221a_1 _11541_ (.A1(_04933_),
    .A2(_04924_),
    .B1(_04932_),
    .B2(_02308_),
    .C1(_05695_),
    .X(_05696_));
 sky130_fd_sc_hd__a21oi_2 _11542_ (.A1(_04853_),
    .A2(_05691_),
    .B1(_05696_),
    .Y(_05697_));
 sky130_fd_sc_hd__nand2_1 _11543_ (.A(_01887_),
    .B(_05676_),
    .Y(_05698_));
 sky130_fd_sc_hd__or2_1 _11544_ (.A(_01887_),
    .B(_05676_),
    .X(_05699_));
 sky130_fd_sc_hd__a22o_1 _11545_ (.A1(\cycles[27] ),
    .A2(_04393_),
    .B1(_04390_),
    .B2(\cycles[59] ),
    .X(_05700_));
 sky130_fd_sc_hd__a221o_1 _11546_ (.A1(\instret[27] ),
    .A2(_04385_),
    .B1(_05072_),
    .B2(\instret[59] ),
    .C1(_05700_),
    .X(_05701_));
 sky130_fd_sc_hd__a221o_1 _11547_ (.A1(_01887_),
    .A2(_05352_),
    .B1(_04376_),
    .B2(_05701_),
    .C1(_01527_),
    .X(_05702_));
 sky130_fd_sc_hd__a31o_1 _11548_ (.A1(_05299_),
    .A2(_05698_),
    .A3(_05699_),
    .B1(_05702_),
    .X(_05703_));
 sky130_fd_sc_hd__a21o_1 _11549_ (.A1(net21),
    .A2(_05033_),
    .B1(_05396_),
    .X(_05704_));
 sky130_fd_sc_hd__a21oi_1 _11550_ (.A1(_04945_),
    .A2(_05704_),
    .B1(_01984_),
    .Y(_05705_));
 sky130_fd_sc_hd__nor2_1 _11551_ (.A(_05032_),
    .B(_05705_),
    .Y(_05706_));
 sky130_fd_sc_hd__o21a_1 _11552_ (.A1(_05697_),
    .A2(_05703_),
    .B1(_05706_),
    .X(_05707_));
 sky130_fd_sc_hd__clkbuf_4 _11553_ (.A(_05707_),
    .X(_05708_));
 sky130_fd_sc_hd__mux2_1 _11554_ (.A0(_05708_),
    .A1(\regs[9][27] ),
    .S(_05515_),
    .X(_05709_));
 sky130_fd_sc_hd__clkbuf_1 _11555_ (.A(_05709_),
    .X(_00346_));
 sky130_fd_sc_hd__xnor2_1 _11556_ (.A(_01917_),
    .B(_05698_),
    .Y(_05710_));
 sky130_fd_sc_hd__a22o_1 _11557_ (.A1(\cycles[28] ),
    .A2(_05073_),
    .B1(_04939_),
    .B2(\cycles[60] ),
    .X(_05711_));
 sky130_fd_sc_hd__a221o_1 _11558_ (.A1(\instret[28] ),
    .A2(_04896_),
    .B1(_05072_),
    .B2(\instret[60] ),
    .C1(_05711_),
    .X(_05712_));
 sky130_fd_sc_hd__a221o_1 _11559_ (.A1(_01917_),
    .A2(_05352_),
    .B1(_04938_),
    .B2(_05712_),
    .C1(_01527_),
    .X(_05713_));
 sky130_fd_sc_hd__nand2_1 _11560_ (.A(_01736_),
    .B(_04587_),
    .Y(_05714_));
 sky130_fd_sc_hd__mux2_1 _11561_ (.A0(_04827_),
    .A1(_04723_),
    .S(_05714_),
    .X(_05715_));
 sky130_fd_sc_hd__nor2_1 _11562_ (.A(_01736_),
    .B(_04587_),
    .Y(_05716_));
 sky130_fd_sc_hd__a21o_1 _11563_ (.A1(_01971_),
    .A2(_05715_),
    .B1(_05716_),
    .X(_05717_));
 sky130_fd_sc_hd__o221a_1 _11564_ (.A1(_04791_),
    .A2(_04881_),
    .B1(_04889_),
    .B2(_04917_),
    .C1(_05717_),
    .X(_05718_));
 sky130_fd_sc_hd__nor2_1 _11565_ (.A(_04571_),
    .B(_04576_),
    .Y(_05719_));
 sky130_fd_sc_hd__o211a_1 _11566_ (.A1(_04561_),
    .A2(_04566_),
    .B1(_05719_),
    .C1(_04562_),
    .X(_05720_));
 sky130_fd_sc_hd__a211o_1 _11567_ (.A1(_04569_),
    .A2(_05693_),
    .B1(_05720_),
    .C1(_05692_),
    .X(_05721_));
 sky130_fd_sc_hd__a31o_1 _11568_ (.A1(_04563_),
    .A2(_05643_),
    .A3(_05719_),
    .B1(_05721_),
    .X(_05722_));
 sky130_fd_sc_hd__xor2_1 _11569_ (.A(_04590_),
    .B(_05722_),
    .X(_05723_));
 sky130_fd_sc_hd__and2_1 _11570_ (.A(\leorv32_alu.input1[27] ),
    .B(_04572_),
    .X(_05724_));
 sky130_fd_sc_hd__a31o_1 _11571_ (.A1(\leorv32_alu.input1[26] ),
    .A2(_04568_),
    .A3(_04573_),
    .B1(_05724_),
    .X(_05725_));
 sky130_fd_sc_hd__a31o_1 _11572_ (.A1(_04577_),
    .A2(_04599_),
    .A3(_05664_),
    .B1(_05725_),
    .X(_05726_));
 sky130_fd_sc_hd__o21ba_1 _11573_ (.A1(_04579_),
    .A2(_05613_),
    .B1_N(_05726_),
    .X(_05727_));
 sky130_fd_sc_hd__xor2_1 _11574_ (.A(_04590_),
    .B(_05727_),
    .X(_05728_));
 sky130_fd_sc_hd__a22o_1 _11575_ (.A1(_04868_),
    .A2(_05723_),
    .B1(_05728_),
    .B2(_05070_),
    .X(_05729_));
 sky130_fd_sc_hd__o2bb2a_1 _11576_ (.A1_N(_04402_),
    .A2_N(_05718_),
    .B1(_04864_),
    .B2(_05729_),
    .X(_05730_));
 sky130_fd_sc_hd__a211o_1 _11577_ (.A1(_05299_),
    .A2(_05710_),
    .B1(_05713_),
    .C1(_05730_),
    .X(_05731_));
 sky130_fd_sc_hd__a21o_1 _11578_ (.A1(net22),
    .A2(_04733_),
    .B1(_05395_),
    .X(_05732_));
 sky130_fd_sc_hd__a21o_1 _11579_ (.A1(_04741_),
    .A2(_05732_),
    .B1(_04815_),
    .X(_05733_));
 sky130_fd_sc_hd__and3_2 _11580_ (.A(_04759_),
    .B(_05731_),
    .C(_05733_),
    .X(_05734_));
 sky130_fd_sc_hd__clkbuf_4 _11581_ (.A(_05734_),
    .X(_05735_));
 sky130_fd_sc_hd__mux2_1 _11582_ (.A0(_05735_),
    .A1(\regs[9][28] ),
    .S(_05515_),
    .X(_05736_));
 sky130_fd_sc_hd__clkbuf_1 _11583_ (.A(_05736_),
    .X(_00347_));
 sky130_fd_sc_hd__o21a_1 _11584_ (.A1(\rs2_content[29] ),
    .A2(_04520_),
    .B1(_04498_),
    .X(_05737_));
 sky130_fd_sc_hd__nand2_1 _11585_ (.A(\leorv32_alu.input1[29] ),
    .B(_05737_),
    .Y(_05738_));
 sky130_fd_sc_hd__nor2_1 _11586_ (.A(\leorv32_alu.input1[29] ),
    .B(_05737_),
    .Y(_05739_));
 sky130_fd_sc_hd__o2bb2a_1 _11587_ (.A1_N(_05277_),
    .A2_N(_04583_),
    .B1(_04933_),
    .B2(_04838_),
    .X(_05740_));
 sky130_fd_sc_hd__o221a_1 _11588_ (.A1(_04827_),
    .A2(_05738_),
    .B1(_05739_),
    .B2(_01972_),
    .C1(_05740_),
    .X(_05741_));
 sky130_fd_sc_hd__a21o_1 _11589_ (.A1(_01823_),
    .A2(_04844_),
    .B1(_02308_),
    .X(_05742_));
 sky130_fd_sc_hd__nand2_1 _11590_ (.A(_04589_),
    .B(_05727_),
    .Y(_05743_));
 sky130_fd_sc_hd__nand2_1 _11591_ (.A(_04588_),
    .B(_05743_),
    .Y(_05744_));
 sky130_fd_sc_hd__nand2_1 _11592_ (.A(_04583_),
    .B(_05744_),
    .Y(_05745_));
 sky130_fd_sc_hd__or2_1 _11593_ (.A(_04583_),
    .B(_05744_),
    .X(_05746_));
 sky130_fd_sc_hd__and2_1 _11594_ (.A(_01736_),
    .B(_04587_),
    .X(_05747_));
 sky130_fd_sc_hd__o21ba_1 _11595_ (.A1(_05747_),
    .A2(_05722_),
    .B1_N(_05716_),
    .X(_05748_));
 sky130_fd_sc_hd__xor2_1 _11596_ (.A(_04583_),
    .B(_05748_),
    .X(_05749_));
 sky130_fd_sc_hd__a32o_1 _11597_ (.A1(_05070_),
    .A2(_05745_),
    .A3(_05746_),
    .B1(_05749_),
    .B2(_04868_),
    .X(_05750_));
 sky130_fd_sc_hd__o2bb2a_1 _11598_ (.A1_N(_05741_),
    .A2_N(_05742_),
    .B1(_05750_),
    .B2(_04864_),
    .X(_05751_));
 sky130_fd_sc_hd__and4_1 _11599_ (.A(_01567_),
    .B(_01917_),
    .C(_01887_),
    .D(_05676_),
    .X(_05752_));
 sky130_fd_sc_hd__inv_2 _11600_ (.A(_05752_),
    .Y(_05753_));
 sky130_fd_sc_hd__a31o_1 _11601_ (.A1(_01917_),
    .A2(_01887_),
    .A3(_05676_),
    .B1(_01567_),
    .X(_05754_));
 sky130_fd_sc_hd__a22o_1 _11602_ (.A1(\cycles[29] ),
    .A2(_04393_),
    .B1(_04390_),
    .B2(\cycles[61] ),
    .X(_05755_));
 sky130_fd_sc_hd__a221o_1 _11603_ (.A1(\instret[29] ),
    .A2(_04385_),
    .B1(_05072_),
    .B2(\instret[61] ),
    .C1(_05755_),
    .X(_05756_));
 sky130_fd_sc_hd__a221o_1 _11604_ (.A1(_01567_),
    .A2(_05352_),
    .B1(_04376_),
    .B2(_05756_),
    .C1(_01527_),
    .X(_05757_));
 sky130_fd_sc_hd__a31o_1 _11605_ (.A1(_05299_),
    .A2(_05753_),
    .A3(_05754_),
    .B1(_05757_),
    .X(_05758_));
 sky130_fd_sc_hd__a21o_1 _11606_ (.A1(net23),
    .A2(_05033_),
    .B1(_05396_),
    .X(_05759_));
 sky130_fd_sc_hd__a21oi_1 _11607_ (.A1(_04945_),
    .A2(_05759_),
    .B1(_01984_),
    .Y(_05760_));
 sky130_fd_sc_hd__nor2_1 _11608_ (.A(_05032_),
    .B(_05760_),
    .Y(_05761_));
 sky130_fd_sc_hd__o21a_1 _11609_ (.A1(_05751_),
    .A2(_05758_),
    .B1(_05761_),
    .X(_05762_));
 sky130_fd_sc_hd__buf_2 _11610_ (.A(_05762_),
    .X(_05763_));
 sky130_fd_sc_hd__mux2_1 _11611_ (.A0(_05763_),
    .A1(\regs[9][29] ),
    .S(_05515_),
    .X(_05764_));
 sky130_fd_sc_hd__clkbuf_1 _11612_ (.A(_05764_),
    .X(_00348_));
 sky130_fd_sc_hd__and2_1 _11613_ (.A(_04583_),
    .B(_04590_),
    .X(_05765_));
 sky130_fd_sc_hd__o21ai_1 _11614_ (.A1(_05739_),
    .A2(_05714_),
    .B1(_05738_),
    .Y(_05766_));
 sky130_fd_sc_hd__a21o_1 _11615_ (.A1(_05722_),
    .A2(_05765_),
    .B1(_05766_),
    .X(_05767_));
 sky130_fd_sc_hd__xnor2_1 _11616_ (.A(_04595_),
    .B(_05767_),
    .Y(_05768_));
 sky130_fd_sc_hd__a21o_1 _11617_ (.A1(_04589_),
    .A2(_05727_),
    .B1(_04604_),
    .X(_05769_));
 sky130_fd_sc_hd__a21oi_1 _11618_ (.A1(_04582_),
    .A2(_05769_),
    .B1(_04595_),
    .Y(_05770_));
 sky130_fd_sc_hd__a31o_1 _11619_ (.A1(_04582_),
    .A2(_04595_),
    .A3(_05769_),
    .B1(_04870_),
    .X(_05771_));
 sky130_fd_sc_hd__o21a_1 _11620_ (.A1(_05770_),
    .A2(_05771_),
    .B1(_04853_),
    .X(_05772_));
 sky130_fd_sc_hd__o21ai_1 _11621_ (.A1(_04782_),
    .A2(_05768_),
    .B1(_05772_),
    .Y(_05773_));
 sky130_fd_sc_hd__mux2_1 _11622_ (.A0(_04723_),
    .A1(_04827_),
    .S(_04594_),
    .X(_05774_));
 sky130_fd_sc_hd__a21o_1 _11623_ (.A1(_01972_),
    .A2(_05774_),
    .B1(_04592_),
    .X(_05775_));
 sky130_fd_sc_hd__o221a_1 _11624_ (.A1(_04917_),
    .A2(_04800_),
    .B1(_04807_),
    .B2(_04933_),
    .C1(_05775_),
    .X(_05776_));
 sky130_fd_sc_hd__nand2_1 _11625_ (.A(_04402_),
    .B(_05776_),
    .Y(_05777_));
 sky130_fd_sc_hd__a22o_1 _11626_ (.A1(\cycles[30] ),
    .A2(_05073_),
    .B1(_04939_),
    .B2(\cycles[62] ),
    .X(_05778_));
 sky130_fd_sc_hd__a221o_1 _11627_ (.A1(\instret[30] ),
    .A2(_04896_),
    .B1(_04395_),
    .B2(\instret[62] ),
    .C1(_05778_),
    .X(_05779_));
 sky130_fd_sc_hd__o21ai_1 _11628_ (.A1(_01602_),
    .A2(_05752_),
    .B1(_04825_),
    .Y(_05780_));
 sky130_fd_sc_hd__a21oi_1 _11629_ (.A1(_01602_),
    .A2(_05752_),
    .B1(_05780_),
    .Y(_05781_));
 sky130_fd_sc_hd__a221o_1 _11630_ (.A1(_01602_),
    .A2(_05352_),
    .B1(_04938_),
    .B2(_05779_),
    .C1(_05781_),
    .X(_05782_));
 sky130_fd_sc_hd__a211o_1 _11631_ (.A1(_05773_),
    .A2(_05777_),
    .B1(_05782_),
    .C1(_01528_),
    .X(_05783_));
 sky130_fd_sc_hd__a21o_1 _11632_ (.A1(net25),
    .A2(_04733_),
    .B1(_05395_),
    .X(_05784_));
 sky130_fd_sc_hd__a21o_1 _11633_ (.A1(_04741_),
    .A2(_05784_),
    .B1(_04815_),
    .X(_05785_));
 sky130_fd_sc_hd__and3_1 _11634_ (.A(_04759_),
    .B(_05783_),
    .C(_05785_),
    .X(_05786_));
 sky130_fd_sc_hd__buf_2 _11635_ (.A(_05786_),
    .X(_05787_));
 sky130_fd_sc_hd__mux2_1 _11636_ (.A0(_05787_),
    .A1(\regs[9][30] ),
    .S(_04768_),
    .X(_05788_));
 sky130_fd_sc_hd__clkbuf_1 _11637_ (.A(_05788_),
    .X(_00349_));
 sky130_fd_sc_hd__nand2_1 _11638_ (.A(_01694_),
    .B(_04593_),
    .Y(_05789_));
 sky130_fd_sc_hd__a211o_1 _11639_ (.A1(_05722_),
    .A2(_05765_),
    .B1(_05766_),
    .C1(_04594_),
    .X(_05790_));
 sky130_fd_sc_hd__a21oi_1 _11640_ (.A1(_05789_),
    .A2(_05790_),
    .B1(_04586_),
    .Y(_05791_));
 sky130_fd_sc_hd__a31o_1 _11641_ (.A1(_04586_),
    .A2(_05789_),
    .A3(_05790_),
    .B1(_04782_),
    .X(_05792_));
 sky130_fd_sc_hd__nor2_1 _11642_ (.A(_05791_),
    .B(_05792_),
    .Y(_05793_));
 sky130_fd_sc_hd__a21oi_1 _11643_ (.A1(\leorv32_alu.input1[30] ),
    .A2(_04593_),
    .B1(_05770_),
    .Y(_05794_));
 sky130_fd_sc_hd__xnor2_1 _11644_ (.A(_04586_),
    .B(_05794_),
    .Y(_05795_));
 sky130_fd_sc_hd__nor2_1 _11645_ (.A(_04870_),
    .B(_05795_),
    .Y(_05796_));
 sky130_fd_sc_hd__o21a_1 _11646_ (.A1(_05793_),
    .A2(_05796_),
    .B1(_04178_),
    .X(_05797_));
 sky130_fd_sc_hd__mux4_1 _11647_ (.A0(_04668_),
    .A1(_04710_),
    .A2(_04711_),
    .A3(_04718_),
    .S0(_04926_),
    .S1(_02307_),
    .X(_05798_));
 sky130_fd_sc_hd__a31o_1 _11648_ (.A1(_01689_),
    .A2(\leorv32_alu.input1[31] ),
    .A3(_04584_),
    .B1(_04610_),
    .X(_05799_));
 sky130_fd_sc_hd__a2bb2o_1 _11649_ (.A1_N(_04619_),
    .A2_N(_05798_),
    .B1(_05799_),
    .B2(_02308_),
    .X(_05800_));
 sky130_fd_sc_hd__a22o_1 _11650_ (.A1(\cycles[31] ),
    .A2(_05073_),
    .B1(_04390_),
    .B2(\cycles[63] ),
    .X(_05801_));
 sky130_fd_sc_hd__a221o_1 _11651_ (.A1(\instret[31] ),
    .A2(_04385_),
    .B1(_05072_),
    .B2(\instret[63] ),
    .C1(_05801_),
    .X(_05802_));
 sky130_fd_sc_hd__a221o_1 _11652_ (.A1(_01539_),
    .A2(_05352_),
    .B1(_04938_),
    .B2(_05802_),
    .C1(_01527_),
    .X(_05803_));
 sky130_fd_sc_hd__a21oi_1 _11653_ (.A1(_01602_),
    .A2(_05752_),
    .B1(_01539_),
    .Y(_05804_));
 sky130_fd_sc_hd__o21ai_1 _11654_ (.A1(_04377_),
    .A2(_05753_),
    .B1(_05299_),
    .Y(_05805_));
 sky130_fd_sc_hd__nor2_1 _11655_ (.A(_05804_),
    .B(_05805_),
    .Y(_05806_));
 sky130_fd_sc_hd__a211o_1 _11656_ (.A1(_04864_),
    .A2(_05800_),
    .B1(_05803_),
    .C1(_05806_),
    .X(_05807_));
 sky130_fd_sc_hd__a21o_1 _11657_ (.A1(net26),
    .A2(_05033_),
    .B1(_05396_),
    .X(_05808_));
 sky130_fd_sc_hd__a21o_1 _11658_ (.A1(_04945_),
    .A2(_05808_),
    .B1(_04949_),
    .X(_05809_));
 sky130_fd_sc_hd__o211a_1 _11659_ (.A1(_05797_),
    .A2(_05807_),
    .B1(_05809_),
    .C1(_04771_),
    .X(_05810_));
 sky130_fd_sc_hd__clkbuf_4 _11660_ (.A(_05810_),
    .X(_05811_));
 sky130_fd_sc_hd__mux2_1 _11661_ (.A0(_05811_),
    .A1(\regs[9][31] ),
    .S(_04768_),
    .X(_05812_));
 sky130_fd_sc_hd__clkbuf_1 _11662_ (.A(_05812_),
    .X(_00350_));
 sky130_fd_sc_hd__clkbuf_4 _11663_ (.A(_04761_),
    .X(_05813_));
 sky130_fd_sc_hd__and3_2 _11664_ (.A(_01648_),
    .B(_01642_),
    .C(_04765_),
    .X(_05814_));
 sky130_fd_sc_hd__and4bb_1 _11665_ (.A_N(_02313_),
    .B_N(_02315_),
    .C(_02241_),
    .D(_04765_),
    .X(_05815_));
 sky130_fd_sc_hd__and2_2 _11666_ (.A(_05814_),
    .B(_05815_),
    .X(_05816_));
 sky130_fd_sc_hd__buf_6 _11667_ (.A(_05816_),
    .X(_05817_));
 sky130_fd_sc_hd__mux2_1 _11668_ (.A0(\regs[7][0] ),
    .A1(_05813_),
    .S(_05817_),
    .X(_05818_));
 sky130_fd_sc_hd__clkbuf_1 _11669_ (.A(_05818_),
    .X(_00351_));
 sky130_fd_sc_hd__clkbuf_4 _11670_ (.A(_04817_),
    .X(_05819_));
 sky130_fd_sc_hd__mux2_1 _11671_ (.A0(\regs[7][1] ),
    .A1(_05819_),
    .S(_05817_),
    .X(_05820_));
 sky130_fd_sc_hd__clkbuf_1 _11672_ (.A(_05820_),
    .X(_00352_));
 sky130_fd_sc_hd__buf_2 _11673_ (.A(_04857_),
    .X(_05821_));
 sky130_fd_sc_hd__mux2_1 _11674_ (.A0(\regs[7][2] ),
    .A1(_05821_),
    .S(_05817_),
    .X(_05822_));
 sky130_fd_sc_hd__clkbuf_1 _11675_ (.A(_05822_),
    .X(_00353_));
 sky130_fd_sc_hd__buf_2 _11676_ (.A(_04903_),
    .X(_05823_));
 sky130_fd_sc_hd__mux2_1 _11677_ (.A0(\regs[7][3] ),
    .A1(_05823_),
    .S(_05817_),
    .X(_05824_));
 sky130_fd_sc_hd__clkbuf_1 _11678_ (.A(_05824_),
    .X(_00354_));
 sky130_fd_sc_hd__buf_2 _11679_ (.A(_04951_),
    .X(_05825_));
 sky130_fd_sc_hd__mux2_1 _11680_ (.A0(\regs[7][4] ),
    .A1(_05825_),
    .S(_05817_),
    .X(_05826_));
 sky130_fd_sc_hd__clkbuf_1 _11681_ (.A(_05826_),
    .X(_00355_));
 sky130_fd_sc_hd__buf_2 _11682_ (.A(_04991_),
    .X(_05827_));
 sky130_fd_sc_hd__mux2_1 _11683_ (.A0(\regs[7][5] ),
    .A1(_05827_),
    .S(_05817_),
    .X(_05828_));
 sky130_fd_sc_hd__clkbuf_1 _11684_ (.A(_05828_),
    .X(_00356_));
 sky130_fd_sc_hd__buf_2 _11685_ (.A(_05029_),
    .X(_05829_));
 sky130_fd_sc_hd__mux2_1 _11686_ (.A0(\regs[7][6] ),
    .A1(_05829_),
    .S(_05817_),
    .X(_05830_));
 sky130_fd_sc_hd__clkbuf_1 _11687_ (.A(_05830_),
    .X(_00357_));
 sky130_fd_sc_hd__buf_2 _11688_ (.A(_05079_),
    .X(_05831_));
 sky130_fd_sc_hd__mux2_1 _11689_ (.A0(\regs[7][7] ),
    .A1(_05831_),
    .S(_05817_),
    .X(_05832_));
 sky130_fd_sc_hd__clkbuf_1 _11690_ (.A(_05832_),
    .X(_00358_));
 sky130_fd_sc_hd__buf_2 _11691_ (.A(_05120_),
    .X(_05833_));
 sky130_fd_sc_hd__mux2_1 _11692_ (.A0(\regs[7][8] ),
    .A1(_05833_),
    .S(_05817_),
    .X(_05834_));
 sky130_fd_sc_hd__clkbuf_1 _11693_ (.A(_05834_),
    .X(_00359_));
 sky130_fd_sc_hd__buf_2 _11694_ (.A(_05156_),
    .X(_05835_));
 sky130_fd_sc_hd__mux2_1 _11695_ (.A0(\regs[7][9] ),
    .A1(_05835_),
    .S(_05817_),
    .X(_05836_));
 sky130_fd_sc_hd__clkbuf_1 _11696_ (.A(_05836_),
    .X(_00360_));
 sky130_fd_sc_hd__clkbuf_4 _11697_ (.A(_05186_),
    .X(_05837_));
 sky130_fd_sc_hd__clkbuf_8 _11698_ (.A(_05816_),
    .X(_05838_));
 sky130_fd_sc_hd__mux2_1 _11699_ (.A0(\regs[7][10] ),
    .A1(_05837_),
    .S(_05838_),
    .X(_05839_));
 sky130_fd_sc_hd__clkbuf_1 _11700_ (.A(_05839_),
    .X(_00361_));
 sky130_fd_sc_hd__clkbuf_4 _11701_ (.A(_05223_),
    .X(_05840_));
 sky130_fd_sc_hd__mux2_1 _11702_ (.A0(\regs[7][11] ),
    .A1(_05840_),
    .S(_05838_),
    .X(_05841_));
 sky130_fd_sc_hd__clkbuf_1 _11703_ (.A(_05841_),
    .X(_00362_));
 sky130_fd_sc_hd__clkbuf_4 _11704_ (.A(_05262_),
    .X(_05842_));
 sky130_fd_sc_hd__mux2_1 _11705_ (.A0(\regs[7][12] ),
    .A1(_05842_),
    .S(_05838_),
    .X(_05843_));
 sky130_fd_sc_hd__clkbuf_1 _11706_ (.A(_05843_),
    .X(_00363_));
 sky130_fd_sc_hd__buf_2 _11707_ (.A(_05295_),
    .X(_05844_));
 sky130_fd_sc_hd__mux2_1 _11708_ (.A0(\regs[7][13] ),
    .A1(_05844_),
    .S(_05838_),
    .X(_05845_));
 sky130_fd_sc_hd__clkbuf_1 _11709_ (.A(_05845_),
    .X(_00364_));
 sky130_fd_sc_hd__clkbuf_4 _11710_ (.A(_05328_),
    .X(_05846_));
 sky130_fd_sc_hd__mux2_1 _11711_ (.A0(\regs[7][14] ),
    .A1(_05846_),
    .S(_05838_),
    .X(_05847_));
 sky130_fd_sc_hd__clkbuf_1 _11712_ (.A(_05847_),
    .X(_00365_));
 sky130_fd_sc_hd__buf_2 _11713_ (.A(_05358_),
    .X(_05848_));
 sky130_fd_sc_hd__mux2_1 _11714_ (.A0(\regs[7][15] ),
    .A1(_05848_),
    .S(_05838_),
    .X(_05849_));
 sky130_fd_sc_hd__clkbuf_1 _11715_ (.A(_05849_),
    .X(_00366_));
 sky130_fd_sc_hd__clkbuf_4 _11716_ (.A(_05399_),
    .X(_05850_));
 sky130_fd_sc_hd__mux2_1 _11717_ (.A0(\regs[7][16] ),
    .A1(_05850_),
    .S(_05838_),
    .X(_05851_));
 sky130_fd_sc_hd__clkbuf_1 _11718_ (.A(_05851_),
    .X(_00367_));
 sky130_fd_sc_hd__clkbuf_4 _11719_ (.A(_05423_),
    .X(_05852_));
 sky130_fd_sc_hd__mux2_1 _11720_ (.A0(\regs[7][17] ),
    .A1(_05852_),
    .S(_05838_),
    .X(_05853_));
 sky130_fd_sc_hd__clkbuf_1 _11721_ (.A(_05853_),
    .X(_00368_));
 sky130_fd_sc_hd__clkbuf_4 _11722_ (.A(_05451_),
    .X(_05854_));
 sky130_fd_sc_hd__mux2_1 _11723_ (.A0(\regs[7][18] ),
    .A1(_05854_),
    .S(_05838_),
    .X(_05855_));
 sky130_fd_sc_hd__clkbuf_1 _11724_ (.A(_05855_),
    .X(_00369_));
 sky130_fd_sc_hd__clkbuf_4 _11725_ (.A(_05476_),
    .X(_05856_));
 sky130_fd_sc_hd__mux2_1 _11726_ (.A0(\regs[7][19] ),
    .A1(_05856_),
    .S(_05838_),
    .X(_05857_));
 sky130_fd_sc_hd__clkbuf_1 _11727_ (.A(_05857_),
    .X(_00370_));
 sky130_fd_sc_hd__buf_2 _11728_ (.A(_05513_),
    .X(_05858_));
 sky130_fd_sc_hd__buf_8 _11729_ (.A(_05816_),
    .X(_05859_));
 sky130_fd_sc_hd__mux2_1 _11730_ (.A0(\regs[7][20] ),
    .A1(_05858_),
    .S(_05859_),
    .X(_05860_));
 sky130_fd_sc_hd__clkbuf_1 _11731_ (.A(_05860_),
    .X(_00371_));
 sky130_fd_sc_hd__clkbuf_4 _11732_ (.A(_05540_),
    .X(_05861_));
 sky130_fd_sc_hd__mux2_1 _11733_ (.A0(\regs[7][21] ),
    .A1(_05861_),
    .S(_05859_),
    .X(_05862_));
 sky130_fd_sc_hd__clkbuf_1 _11734_ (.A(_05862_),
    .X(_00372_));
 sky130_fd_sc_hd__clkbuf_4 _11735_ (.A(_05569_),
    .X(_05863_));
 sky130_fd_sc_hd__mux2_1 _11736_ (.A0(\regs[7][22] ),
    .A1(_05863_),
    .S(_05859_),
    .X(_05864_));
 sky130_fd_sc_hd__clkbuf_1 _11737_ (.A(_05864_),
    .X(_00373_));
 sky130_fd_sc_hd__buf_2 _11738_ (.A(_05599_),
    .X(_05865_));
 sky130_fd_sc_hd__mux2_1 _11739_ (.A0(\regs[7][23] ),
    .A1(_05865_),
    .S(_05859_),
    .X(_05866_));
 sky130_fd_sc_hd__clkbuf_1 _11740_ (.A(_05866_),
    .X(_00374_));
 sky130_fd_sc_hd__clkbuf_4 _11741_ (.A(_05635_),
    .X(_05867_));
 sky130_fd_sc_hd__mux2_1 _11742_ (.A0(\regs[7][24] ),
    .A1(_05867_),
    .S(_05859_),
    .X(_05868_));
 sky130_fd_sc_hd__clkbuf_1 _11743_ (.A(_05868_),
    .X(_00375_));
 sky130_fd_sc_hd__buf_2 _11744_ (.A(_05659_),
    .X(_05869_));
 sky130_fd_sc_hd__mux2_1 _11745_ (.A0(\regs[7][25] ),
    .A1(_05869_),
    .S(_05859_),
    .X(_05870_));
 sky130_fd_sc_hd__clkbuf_1 _11746_ (.A(_05870_),
    .X(_00376_));
 sky130_fd_sc_hd__clkbuf_4 _11747_ (.A(_05683_),
    .X(_05871_));
 sky130_fd_sc_hd__mux2_1 _11748_ (.A0(\regs[7][26] ),
    .A1(_05871_),
    .S(_05859_),
    .X(_05872_));
 sky130_fd_sc_hd__clkbuf_1 _11749_ (.A(_05872_),
    .X(_00377_));
 sky130_fd_sc_hd__clkbuf_4 _11750_ (.A(_05707_),
    .X(_05873_));
 sky130_fd_sc_hd__mux2_1 _11751_ (.A0(\regs[7][27] ),
    .A1(_05873_),
    .S(_05859_),
    .X(_05874_));
 sky130_fd_sc_hd__clkbuf_1 _11752_ (.A(_05874_),
    .X(_00378_));
 sky130_fd_sc_hd__buf_2 _11753_ (.A(_05734_),
    .X(_05875_));
 sky130_fd_sc_hd__mux2_1 _11754_ (.A0(\regs[7][28] ),
    .A1(_05875_),
    .S(_05859_),
    .X(_05876_));
 sky130_fd_sc_hd__clkbuf_1 _11755_ (.A(_05876_),
    .X(_00379_));
 sky130_fd_sc_hd__clkbuf_4 _11756_ (.A(_05762_),
    .X(_05877_));
 sky130_fd_sc_hd__mux2_1 _11757_ (.A0(\regs[7][29] ),
    .A1(_05877_),
    .S(_05859_),
    .X(_05878_));
 sky130_fd_sc_hd__clkbuf_1 _11758_ (.A(_05878_),
    .X(_00380_));
 sky130_fd_sc_hd__buf_2 _11759_ (.A(_05786_),
    .X(_05879_));
 sky130_fd_sc_hd__mux2_1 _11760_ (.A0(\regs[7][30] ),
    .A1(_05879_),
    .S(_05816_),
    .X(_05880_));
 sky130_fd_sc_hd__clkbuf_1 _11761_ (.A(_05880_),
    .X(_00381_));
 sky130_fd_sc_hd__buf_2 _11762_ (.A(_05810_),
    .X(_05881_));
 sky130_fd_sc_hd__mux2_1 _11763_ (.A0(\regs[7][31] ),
    .A1(_05881_),
    .S(_05816_),
    .X(_05882_));
 sky130_fd_sc_hd__clkbuf_1 _11764_ (.A(_05882_),
    .X(_00382_));
 sky130_fd_sc_hd__nand3b_4 _11765_ (.A_N(_01642_),
    .B(_04756_),
    .C(_01648_),
    .Y(_05883_));
 sky130_fd_sc_hd__inv_2 _11766_ (.A(_05883_),
    .Y(_05884_));
 sky130_fd_sc_hd__nand2_4 _11767_ (.A(_04767_),
    .B(_05884_),
    .Y(_05885_));
 sky130_fd_sc_hd__clkbuf_8 _11768_ (.A(_05885_),
    .X(_05886_));
 sky130_fd_sc_hd__mux2_1 _11769_ (.A0(_04762_),
    .A1(\regs[10][0] ),
    .S(_05886_),
    .X(_05887_));
 sky130_fd_sc_hd__clkbuf_1 _11770_ (.A(_05887_),
    .X(_00383_));
 sky130_fd_sc_hd__mux2_1 _11771_ (.A0(_04818_),
    .A1(\regs[10][1] ),
    .S(_05886_),
    .X(_05888_));
 sky130_fd_sc_hd__clkbuf_1 _11772_ (.A(_05888_),
    .X(_00384_));
 sky130_fd_sc_hd__mux2_1 _11773_ (.A0(_04858_),
    .A1(\regs[10][2] ),
    .S(_05886_),
    .X(_05889_));
 sky130_fd_sc_hd__clkbuf_1 _11774_ (.A(_05889_),
    .X(_00385_));
 sky130_fd_sc_hd__mux2_1 _11775_ (.A0(_04904_),
    .A1(\regs[10][3] ),
    .S(_05886_),
    .X(_05890_));
 sky130_fd_sc_hd__clkbuf_1 _11776_ (.A(_05890_),
    .X(_00386_));
 sky130_fd_sc_hd__mux2_1 _11777_ (.A0(_04952_),
    .A1(\regs[10][4] ),
    .S(_05886_),
    .X(_05891_));
 sky130_fd_sc_hd__clkbuf_1 _11778_ (.A(_05891_),
    .X(_00387_));
 sky130_fd_sc_hd__mux2_1 _11779_ (.A0(_04992_),
    .A1(\regs[10][5] ),
    .S(_05886_),
    .X(_05892_));
 sky130_fd_sc_hd__clkbuf_1 _11780_ (.A(_05892_),
    .X(_00388_));
 sky130_fd_sc_hd__mux2_1 _11781_ (.A0(_05030_),
    .A1(\regs[10][6] ),
    .S(_05886_),
    .X(_05893_));
 sky130_fd_sc_hd__clkbuf_1 _11782_ (.A(_05893_),
    .X(_00389_));
 sky130_fd_sc_hd__mux2_1 _11783_ (.A0(_05080_),
    .A1(\regs[10][7] ),
    .S(_05886_),
    .X(_05894_));
 sky130_fd_sc_hd__clkbuf_1 _11784_ (.A(_05894_),
    .X(_00390_));
 sky130_fd_sc_hd__mux2_1 _11785_ (.A0(_05121_),
    .A1(\regs[10][8] ),
    .S(_05886_),
    .X(_05895_));
 sky130_fd_sc_hd__clkbuf_1 _11786_ (.A(_05895_),
    .X(_00391_));
 sky130_fd_sc_hd__mux2_1 _11787_ (.A0(_05157_),
    .A1(\regs[10][9] ),
    .S(_05886_),
    .X(_05896_));
 sky130_fd_sc_hd__clkbuf_1 _11788_ (.A(_05896_),
    .X(_00392_));
 sky130_fd_sc_hd__buf_4 _11789_ (.A(_05885_),
    .X(_05897_));
 sky130_fd_sc_hd__mux2_1 _11790_ (.A0(_05187_),
    .A1(\regs[10][10] ),
    .S(_05897_),
    .X(_05898_));
 sky130_fd_sc_hd__clkbuf_1 _11791_ (.A(_05898_),
    .X(_00393_));
 sky130_fd_sc_hd__mux2_1 _11792_ (.A0(_05224_),
    .A1(\regs[10][11] ),
    .S(_05897_),
    .X(_05899_));
 sky130_fd_sc_hd__clkbuf_1 _11793_ (.A(_05899_),
    .X(_00394_));
 sky130_fd_sc_hd__mux2_1 _11794_ (.A0(_05263_),
    .A1(\regs[10][12] ),
    .S(_05897_),
    .X(_05900_));
 sky130_fd_sc_hd__clkbuf_1 _11795_ (.A(_05900_),
    .X(_00395_));
 sky130_fd_sc_hd__mux2_1 _11796_ (.A0(_05296_),
    .A1(\regs[10][13] ),
    .S(_05897_),
    .X(_05901_));
 sky130_fd_sc_hd__clkbuf_1 _11797_ (.A(_05901_),
    .X(_00396_));
 sky130_fd_sc_hd__mux2_1 _11798_ (.A0(_05329_),
    .A1(\regs[10][14] ),
    .S(_05897_),
    .X(_05902_));
 sky130_fd_sc_hd__clkbuf_1 _11799_ (.A(_05902_),
    .X(_00397_));
 sky130_fd_sc_hd__mux2_1 _11800_ (.A0(_05359_),
    .A1(\regs[10][15] ),
    .S(_05897_),
    .X(_05903_));
 sky130_fd_sc_hd__clkbuf_1 _11801_ (.A(_05903_),
    .X(_00398_));
 sky130_fd_sc_hd__mux2_1 _11802_ (.A0(_05400_),
    .A1(\regs[10][16] ),
    .S(_05897_),
    .X(_05904_));
 sky130_fd_sc_hd__clkbuf_1 _11803_ (.A(_05904_),
    .X(_00399_));
 sky130_fd_sc_hd__mux2_1 _11804_ (.A0(_05424_),
    .A1(\regs[10][17] ),
    .S(_05897_),
    .X(_05905_));
 sky130_fd_sc_hd__clkbuf_1 _11805_ (.A(_05905_),
    .X(_00400_));
 sky130_fd_sc_hd__mux2_1 _11806_ (.A0(_05452_),
    .A1(\regs[10][18] ),
    .S(_05897_),
    .X(_05906_));
 sky130_fd_sc_hd__clkbuf_1 _11807_ (.A(_05906_),
    .X(_00401_));
 sky130_fd_sc_hd__mux2_1 _11808_ (.A0(_05477_),
    .A1(\regs[10][19] ),
    .S(_05897_),
    .X(_05907_));
 sky130_fd_sc_hd__clkbuf_1 _11809_ (.A(_05907_),
    .X(_00402_));
 sky130_fd_sc_hd__buf_8 _11810_ (.A(_05885_),
    .X(_05908_));
 sky130_fd_sc_hd__mux2_1 _11811_ (.A0(_05514_),
    .A1(\regs[10][20] ),
    .S(_05908_),
    .X(_05909_));
 sky130_fd_sc_hd__clkbuf_1 _11812_ (.A(_05909_),
    .X(_00403_));
 sky130_fd_sc_hd__mux2_1 _11813_ (.A0(_05541_),
    .A1(\regs[10][21] ),
    .S(_05908_),
    .X(_05910_));
 sky130_fd_sc_hd__clkbuf_1 _11814_ (.A(_05910_),
    .X(_00404_));
 sky130_fd_sc_hd__mux2_1 _11815_ (.A0(_05570_),
    .A1(\regs[10][22] ),
    .S(_05908_),
    .X(_05911_));
 sky130_fd_sc_hd__clkbuf_1 _11816_ (.A(_05911_),
    .X(_00405_));
 sky130_fd_sc_hd__mux2_1 _11817_ (.A0(_05600_),
    .A1(\regs[10][23] ),
    .S(_05908_),
    .X(_05912_));
 sky130_fd_sc_hd__clkbuf_1 _11818_ (.A(_05912_),
    .X(_00406_));
 sky130_fd_sc_hd__mux2_1 _11819_ (.A0(_05636_),
    .A1(\regs[10][24] ),
    .S(_05908_),
    .X(_05913_));
 sky130_fd_sc_hd__clkbuf_1 _11820_ (.A(_05913_),
    .X(_00407_));
 sky130_fd_sc_hd__mux2_1 _11821_ (.A0(_05660_),
    .A1(\regs[10][25] ),
    .S(_05908_),
    .X(_05914_));
 sky130_fd_sc_hd__clkbuf_1 _11822_ (.A(_05914_),
    .X(_00408_));
 sky130_fd_sc_hd__mux2_1 _11823_ (.A0(_05684_),
    .A1(\regs[10][26] ),
    .S(_05908_),
    .X(_05915_));
 sky130_fd_sc_hd__clkbuf_1 _11824_ (.A(_05915_),
    .X(_00409_));
 sky130_fd_sc_hd__mux2_1 _11825_ (.A0(_05708_),
    .A1(\regs[10][27] ),
    .S(_05908_),
    .X(_05916_));
 sky130_fd_sc_hd__clkbuf_1 _11826_ (.A(_05916_),
    .X(_00410_));
 sky130_fd_sc_hd__mux2_1 _11827_ (.A0(_05735_),
    .A1(\regs[10][28] ),
    .S(_05908_),
    .X(_05917_));
 sky130_fd_sc_hd__clkbuf_1 _11828_ (.A(_05917_),
    .X(_00411_));
 sky130_fd_sc_hd__mux2_1 _11829_ (.A0(_05763_),
    .A1(\regs[10][29] ),
    .S(_05908_),
    .X(_05918_));
 sky130_fd_sc_hd__clkbuf_1 _11830_ (.A(_05918_),
    .X(_00412_));
 sky130_fd_sc_hd__mux2_1 _11831_ (.A0(_05787_),
    .A1(\regs[10][30] ),
    .S(_05885_),
    .X(_05919_));
 sky130_fd_sc_hd__clkbuf_1 _11832_ (.A(_05919_),
    .X(_00413_));
 sky130_fd_sc_hd__mux2_1 _11833_ (.A0(_05811_),
    .A1(\regs[10][31] ),
    .S(_05885_),
    .X(_05920_));
 sky130_fd_sc_hd__clkbuf_1 _11834_ (.A(_05920_),
    .X(_00414_));
 sky130_fd_sc_hd__or3b_4 _11835_ (.A(_04766_),
    .B(_02313_),
    .C_N(_02241_),
    .X(_05921_));
 sky130_fd_sc_hd__nor2_4 _11836_ (.A(_04758_),
    .B(_05921_),
    .Y(_05922_));
 sky130_fd_sc_hd__clkbuf_8 _11837_ (.A(_05922_),
    .X(_05923_));
 sky130_fd_sc_hd__mux2_1 _11838_ (.A0(\regs[12][0] ),
    .A1(_05813_),
    .S(_05923_),
    .X(_05924_));
 sky130_fd_sc_hd__clkbuf_1 _11839_ (.A(_05924_),
    .X(_00415_));
 sky130_fd_sc_hd__mux2_1 _11840_ (.A0(\regs[12][1] ),
    .A1(_05819_),
    .S(_05923_),
    .X(_05925_));
 sky130_fd_sc_hd__clkbuf_1 _11841_ (.A(_05925_),
    .X(_00416_));
 sky130_fd_sc_hd__mux2_1 _11842_ (.A0(\regs[12][2] ),
    .A1(_05821_),
    .S(_05923_),
    .X(_05926_));
 sky130_fd_sc_hd__clkbuf_1 _11843_ (.A(_05926_),
    .X(_00417_));
 sky130_fd_sc_hd__mux2_1 _11844_ (.A0(\regs[12][3] ),
    .A1(_05823_),
    .S(_05923_),
    .X(_05927_));
 sky130_fd_sc_hd__clkbuf_1 _11845_ (.A(_05927_),
    .X(_00418_));
 sky130_fd_sc_hd__mux2_1 _11846_ (.A0(\regs[12][4] ),
    .A1(_05825_),
    .S(_05923_),
    .X(_05928_));
 sky130_fd_sc_hd__clkbuf_1 _11847_ (.A(_05928_),
    .X(_00419_));
 sky130_fd_sc_hd__mux2_1 _11848_ (.A0(\regs[12][5] ),
    .A1(_05827_),
    .S(_05923_),
    .X(_05929_));
 sky130_fd_sc_hd__clkbuf_1 _11849_ (.A(_05929_),
    .X(_00420_));
 sky130_fd_sc_hd__mux2_1 _11850_ (.A0(\regs[12][6] ),
    .A1(_05829_),
    .S(_05923_),
    .X(_05930_));
 sky130_fd_sc_hd__clkbuf_1 _11851_ (.A(_05930_),
    .X(_00421_));
 sky130_fd_sc_hd__mux2_1 _11852_ (.A0(\regs[12][7] ),
    .A1(_05831_),
    .S(_05923_),
    .X(_05931_));
 sky130_fd_sc_hd__clkbuf_1 _11853_ (.A(_05931_),
    .X(_00422_));
 sky130_fd_sc_hd__mux2_1 _11854_ (.A0(\regs[12][8] ),
    .A1(_05833_),
    .S(_05923_),
    .X(_05932_));
 sky130_fd_sc_hd__clkbuf_1 _11855_ (.A(_05932_),
    .X(_00423_));
 sky130_fd_sc_hd__mux2_1 _11856_ (.A0(\regs[12][9] ),
    .A1(_05835_),
    .S(_05923_),
    .X(_05933_));
 sky130_fd_sc_hd__clkbuf_1 _11857_ (.A(_05933_),
    .X(_00424_));
 sky130_fd_sc_hd__clkbuf_8 _11858_ (.A(_05922_),
    .X(_05934_));
 sky130_fd_sc_hd__mux2_1 _11859_ (.A0(\regs[12][10] ),
    .A1(_05837_),
    .S(_05934_),
    .X(_05935_));
 sky130_fd_sc_hd__clkbuf_1 _11860_ (.A(_05935_),
    .X(_00425_));
 sky130_fd_sc_hd__mux2_1 _11861_ (.A0(\regs[12][11] ),
    .A1(_05840_),
    .S(_05934_),
    .X(_05936_));
 sky130_fd_sc_hd__clkbuf_1 _11862_ (.A(_05936_),
    .X(_00426_));
 sky130_fd_sc_hd__mux2_1 _11863_ (.A0(\regs[12][12] ),
    .A1(_05842_),
    .S(_05934_),
    .X(_05937_));
 sky130_fd_sc_hd__clkbuf_1 _11864_ (.A(_05937_),
    .X(_00427_));
 sky130_fd_sc_hd__mux2_1 _11865_ (.A0(\regs[12][13] ),
    .A1(_05844_),
    .S(_05934_),
    .X(_05938_));
 sky130_fd_sc_hd__clkbuf_1 _11866_ (.A(_05938_),
    .X(_00428_));
 sky130_fd_sc_hd__mux2_1 _11867_ (.A0(\regs[12][14] ),
    .A1(_05846_),
    .S(_05934_),
    .X(_05939_));
 sky130_fd_sc_hd__clkbuf_1 _11868_ (.A(_05939_),
    .X(_00429_));
 sky130_fd_sc_hd__mux2_1 _11869_ (.A0(\regs[12][15] ),
    .A1(_05848_),
    .S(_05934_),
    .X(_05940_));
 sky130_fd_sc_hd__clkbuf_1 _11870_ (.A(_05940_),
    .X(_00430_));
 sky130_fd_sc_hd__mux2_1 _11871_ (.A0(\regs[12][16] ),
    .A1(_05850_),
    .S(_05934_),
    .X(_05941_));
 sky130_fd_sc_hd__clkbuf_1 _11872_ (.A(_05941_),
    .X(_00431_));
 sky130_fd_sc_hd__mux2_1 _11873_ (.A0(\regs[12][17] ),
    .A1(_05852_),
    .S(_05934_),
    .X(_05942_));
 sky130_fd_sc_hd__clkbuf_1 _11874_ (.A(_05942_),
    .X(_00432_));
 sky130_fd_sc_hd__mux2_1 _11875_ (.A0(\regs[12][18] ),
    .A1(_05854_),
    .S(_05934_),
    .X(_05943_));
 sky130_fd_sc_hd__clkbuf_1 _11876_ (.A(_05943_),
    .X(_00433_));
 sky130_fd_sc_hd__mux2_1 _11877_ (.A0(\regs[12][19] ),
    .A1(_05856_),
    .S(_05934_),
    .X(_05944_));
 sky130_fd_sc_hd__clkbuf_1 _11878_ (.A(_05944_),
    .X(_00434_));
 sky130_fd_sc_hd__buf_6 _11879_ (.A(_05922_),
    .X(_05945_));
 sky130_fd_sc_hd__mux2_1 _11880_ (.A0(\regs[12][20] ),
    .A1(_05858_),
    .S(_05945_),
    .X(_05946_));
 sky130_fd_sc_hd__clkbuf_1 _11881_ (.A(_05946_),
    .X(_00435_));
 sky130_fd_sc_hd__mux2_1 _11882_ (.A0(\regs[12][21] ),
    .A1(_05861_),
    .S(_05945_),
    .X(_05947_));
 sky130_fd_sc_hd__clkbuf_1 _11883_ (.A(_05947_),
    .X(_00436_));
 sky130_fd_sc_hd__mux2_1 _11884_ (.A0(\regs[12][22] ),
    .A1(_05863_),
    .S(_05945_),
    .X(_05948_));
 sky130_fd_sc_hd__clkbuf_1 _11885_ (.A(_05948_),
    .X(_00437_));
 sky130_fd_sc_hd__mux2_1 _11886_ (.A0(\regs[12][23] ),
    .A1(_05865_),
    .S(_05945_),
    .X(_05949_));
 sky130_fd_sc_hd__clkbuf_1 _11887_ (.A(_05949_),
    .X(_00438_));
 sky130_fd_sc_hd__mux2_1 _11888_ (.A0(\regs[12][24] ),
    .A1(_05867_),
    .S(_05945_),
    .X(_05950_));
 sky130_fd_sc_hd__clkbuf_1 _11889_ (.A(_05950_),
    .X(_00439_));
 sky130_fd_sc_hd__mux2_1 _11890_ (.A0(\regs[12][25] ),
    .A1(_05869_),
    .S(_05945_),
    .X(_05951_));
 sky130_fd_sc_hd__clkbuf_1 _11891_ (.A(_05951_),
    .X(_00440_));
 sky130_fd_sc_hd__mux2_1 _11892_ (.A0(\regs[12][26] ),
    .A1(_05871_),
    .S(_05945_),
    .X(_05952_));
 sky130_fd_sc_hd__clkbuf_1 _11893_ (.A(_05952_),
    .X(_00441_));
 sky130_fd_sc_hd__mux2_1 _11894_ (.A0(\regs[12][27] ),
    .A1(_05873_),
    .S(_05945_),
    .X(_05953_));
 sky130_fd_sc_hd__clkbuf_1 _11895_ (.A(_05953_),
    .X(_00442_));
 sky130_fd_sc_hd__mux2_1 _11896_ (.A0(\regs[12][28] ),
    .A1(_05875_),
    .S(_05945_),
    .X(_05954_));
 sky130_fd_sc_hd__clkbuf_1 _11897_ (.A(_05954_),
    .X(_00443_));
 sky130_fd_sc_hd__mux2_1 _11898_ (.A0(\regs[12][29] ),
    .A1(_05877_),
    .S(_05945_),
    .X(_05955_));
 sky130_fd_sc_hd__clkbuf_1 _11899_ (.A(_05955_),
    .X(_00444_));
 sky130_fd_sc_hd__mux2_1 _11900_ (.A0(\regs[12][30] ),
    .A1(_05879_),
    .S(_05922_),
    .X(_05956_));
 sky130_fd_sc_hd__clkbuf_1 _11901_ (.A(_05956_),
    .X(_00445_));
 sky130_fd_sc_hd__mux2_1 _11902_ (.A0(\regs[12][31] ),
    .A1(_05881_),
    .S(_05922_),
    .X(_05957_));
 sky130_fd_sc_hd__clkbuf_1 _11903_ (.A(_05957_),
    .X(_00446_));
 sky130_fd_sc_hd__nand3_4 _11904_ (.A(_01648_),
    .B(_01642_),
    .C(_04765_),
    .Y(_05958_));
 sky130_fd_sc_hd__nor2_4 _11905_ (.A(_05958_),
    .B(_05921_),
    .Y(_05959_));
 sky130_fd_sc_hd__clkbuf_8 _11906_ (.A(_05959_),
    .X(_05960_));
 sky130_fd_sc_hd__mux2_1 _11907_ (.A0(\regs[15][0] ),
    .A1(_05813_),
    .S(_05960_),
    .X(_05961_));
 sky130_fd_sc_hd__clkbuf_1 _11908_ (.A(_05961_),
    .X(_00447_));
 sky130_fd_sc_hd__mux2_1 _11909_ (.A0(\regs[15][1] ),
    .A1(_05819_),
    .S(_05960_),
    .X(_05962_));
 sky130_fd_sc_hd__clkbuf_1 _11910_ (.A(_05962_),
    .X(_00448_));
 sky130_fd_sc_hd__mux2_1 _11911_ (.A0(\regs[15][2] ),
    .A1(_05821_),
    .S(_05960_),
    .X(_05963_));
 sky130_fd_sc_hd__clkbuf_1 _11912_ (.A(_05963_),
    .X(_00449_));
 sky130_fd_sc_hd__mux2_1 _11913_ (.A0(\regs[15][3] ),
    .A1(_05823_),
    .S(_05960_),
    .X(_05964_));
 sky130_fd_sc_hd__clkbuf_1 _11914_ (.A(_05964_),
    .X(_00450_));
 sky130_fd_sc_hd__mux2_1 _11915_ (.A0(\regs[15][4] ),
    .A1(_05825_),
    .S(_05960_),
    .X(_05965_));
 sky130_fd_sc_hd__clkbuf_1 _11916_ (.A(_05965_),
    .X(_00451_));
 sky130_fd_sc_hd__mux2_1 _11917_ (.A0(\regs[15][5] ),
    .A1(_05827_),
    .S(_05960_),
    .X(_05966_));
 sky130_fd_sc_hd__clkbuf_1 _11918_ (.A(_05966_),
    .X(_00452_));
 sky130_fd_sc_hd__mux2_1 _11919_ (.A0(\regs[15][6] ),
    .A1(_05829_),
    .S(_05960_),
    .X(_05967_));
 sky130_fd_sc_hd__clkbuf_1 _11920_ (.A(_05967_),
    .X(_00453_));
 sky130_fd_sc_hd__mux2_1 _11921_ (.A0(\regs[15][7] ),
    .A1(_05831_),
    .S(_05960_),
    .X(_05968_));
 sky130_fd_sc_hd__clkbuf_1 _11922_ (.A(_05968_),
    .X(_00454_));
 sky130_fd_sc_hd__mux2_1 _11923_ (.A0(\regs[15][8] ),
    .A1(_05833_),
    .S(_05960_),
    .X(_05969_));
 sky130_fd_sc_hd__clkbuf_1 _11924_ (.A(_05969_),
    .X(_00455_));
 sky130_fd_sc_hd__mux2_1 _11925_ (.A0(\regs[15][9] ),
    .A1(_05835_),
    .S(_05960_),
    .X(_05970_));
 sky130_fd_sc_hd__clkbuf_1 _11926_ (.A(_05970_),
    .X(_00456_));
 sky130_fd_sc_hd__buf_4 _11927_ (.A(_05959_),
    .X(_05971_));
 sky130_fd_sc_hd__mux2_1 _11928_ (.A0(\regs[15][10] ),
    .A1(_05837_),
    .S(_05971_),
    .X(_05972_));
 sky130_fd_sc_hd__clkbuf_1 _11929_ (.A(_05972_),
    .X(_00457_));
 sky130_fd_sc_hd__mux2_1 _11930_ (.A0(\regs[15][11] ),
    .A1(_05840_),
    .S(_05971_),
    .X(_05973_));
 sky130_fd_sc_hd__clkbuf_1 _11931_ (.A(_05973_),
    .X(_00458_));
 sky130_fd_sc_hd__mux2_1 _11932_ (.A0(\regs[15][12] ),
    .A1(_05842_),
    .S(_05971_),
    .X(_05974_));
 sky130_fd_sc_hd__clkbuf_1 _11933_ (.A(_05974_),
    .X(_00459_));
 sky130_fd_sc_hd__mux2_1 _11934_ (.A0(\regs[15][13] ),
    .A1(_05844_),
    .S(_05971_),
    .X(_05975_));
 sky130_fd_sc_hd__clkbuf_1 _11935_ (.A(_05975_),
    .X(_00460_));
 sky130_fd_sc_hd__mux2_1 _11936_ (.A0(\regs[15][14] ),
    .A1(_05846_),
    .S(_05971_),
    .X(_05976_));
 sky130_fd_sc_hd__clkbuf_1 _11937_ (.A(_05976_),
    .X(_00461_));
 sky130_fd_sc_hd__mux2_1 _11938_ (.A0(\regs[15][15] ),
    .A1(_05848_),
    .S(_05971_),
    .X(_05977_));
 sky130_fd_sc_hd__clkbuf_1 _11939_ (.A(_05977_),
    .X(_00462_));
 sky130_fd_sc_hd__mux2_1 _11940_ (.A0(\regs[15][16] ),
    .A1(_05850_),
    .S(_05971_),
    .X(_05978_));
 sky130_fd_sc_hd__clkbuf_1 _11941_ (.A(_05978_),
    .X(_00463_));
 sky130_fd_sc_hd__mux2_1 _11942_ (.A0(\regs[15][17] ),
    .A1(_05852_),
    .S(_05971_),
    .X(_05979_));
 sky130_fd_sc_hd__clkbuf_1 _11943_ (.A(_05979_),
    .X(_00464_));
 sky130_fd_sc_hd__mux2_1 _11944_ (.A0(\regs[15][18] ),
    .A1(_05854_),
    .S(_05971_),
    .X(_05980_));
 sky130_fd_sc_hd__clkbuf_1 _11945_ (.A(_05980_),
    .X(_00465_));
 sky130_fd_sc_hd__mux2_1 _11946_ (.A0(\regs[15][19] ),
    .A1(_05856_),
    .S(_05971_),
    .X(_05981_));
 sky130_fd_sc_hd__clkbuf_1 _11947_ (.A(_05981_),
    .X(_00466_));
 sky130_fd_sc_hd__buf_6 _11948_ (.A(_05959_),
    .X(_05982_));
 sky130_fd_sc_hd__mux2_1 _11949_ (.A0(\regs[15][20] ),
    .A1(_05858_),
    .S(_05982_),
    .X(_05983_));
 sky130_fd_sc_hd__clkbuf_1 _11950_ (.A(_05983_),
    .X(_00467_));
 sky130_fd_sc_hd__mux2_1 _11951_ (.A0(\regs[15][21] ),
    .A1(_05861_),
    .S(_05982_),
    .X(_05984_));
 sky130_fd_sc_hd__clkbuf_1 _11952_ (.A(_05984_),
    .X(_00468_));
 sky130_fd_sc_hd__mux2_1 _11953_ (.A0(\regs[15][22] ),
    .A1(_05863_),
    .S(_05982_),
    .X(_05985_));
 sky130_fd_sc_hd__clkbuf_1 _11954_ (.A(_05985_),
    .X(_00469_));
 sky130_fd_sc_hd__mux2_1 _11955_ (.A0(\regs[15][23] ),
    .A1(_05865_),
    .S(_05982_),
    .X(_05986_));
 sky130_fd_sc_hd__clkbuf_1 _11956_ (.A(_05986_),
    .X(_00470_));
 sky130_fd_sc_hd__mux2_1 _11957_ (.A0(\regs[15][24] ),
    .A1(_05867_),
    .S(_05982_),
    .X(_05987_));
 sky130_fd_sc_hd__clkbuf_1 _11958_ (.A(_05987_),
    .X(_00471_));
 sky130_fd_sc_hd__mux2_1 _11959_ (.A0(\regs[15][25] ),
    .A1(_05869_),
    .S(_05982_),
    .X(_05988_));
 sky130_fd_sc_hd__clkbuf_1 _11960_ (.A(_05988_),
    .X(_00472_));
 sky130_fd_sc_hd__mux2_1 _11961_ (.A0(\regs[15][26] ),
    .A1(_05871_),
    .S(_05982_),
    .X(_05989_));
 sky130_fd_sc_hd__clkbuf_1 _11962_ (.A(_05989_),
    .X(_00473_));
 sky130_fd_sc_hd__mux2_1 _11963_ (.A0(\regs[15][27] ),
    .A1(_05873_),
    .S(_05982_),
    .X(_05990_));
 sky130_fd_sc_hd__clkbuf_1 _11964_ (.A(_05990_),
    .X(_00474_));
 sky130_fd_sc_hd__mux2_1 _11965_ (.A0(\regs[15][28] ),
    .A1(_05875_),
    .S(_05982_),
    .X(_05991_));
 sky130_fd_sc_hd__clkbuf_1 _11966_ (.A(_05991_),
    .X(_00475_));
 sky130_fd_sc_hd__mux2_1 _11967_ (.A0(\regs[15][29] ),
    .A1(_05877_),
    .S(_05982_),
    .X(_05992_));
 sky130_fd_sc_hd__clkbuf_1 _11968_ (.A(_05992_),
    .X(_00476_));
 sky130_fd_sc_hd__mux2_1 _11969_ (.A0(\regs[15][30] ),
    .A1(_05879_),
    .S(_05959_),
    .X(_05993_));
 sky130_fd_sc_hd__clkbuf_1 _11970_ (.A(_05993_),
    .X(_00477_));
 sky130_fd_sc_hd__mux2_1 _11971_ (.A0(\regs[15][31] ),
    .A1(_05881_),
    .S(_05959_),
    .X(_05994_));
 sky130_fd_sc_hd__clkbuf_1 _11972_ (.A(_05994_),
    .X(_00478_));
 sky130_fd_sc_hd__and2_4 _11973_ (.A(_04764_),
    .B(_05815_),
    .X(_05995_));
 sky130_fd_sc_hd__buf_6 _11974_ (.A(_05995_),
    .X(_05996_));
 sky130_fd_sc_hd__mux2_1 _11975_ (.A0(\regs[5][0] ),
    .A1(_05813_),
    .S(_05996_),
    .X(_05997_));
 sky130_fd_sc_hd__clkbuf_1 _11976_ (.A(_05997_),
    .X(_00479_));
 sky130_fd_sc_hd__mux2_1 _11977_ (.A0(\regs[5][1] ),
    .A1(_05819_),
    .S(_05996_),
    .X(_05998_));
 sky130_fd_sc_hd__clkbuf_1 _11978_ (.A(_05998_),
    .X(_00480_));
 sky130_fd_sc_hd__mux2_1 _11979_ (.A0(\regs[5][2] ),
    .A1(_05821_),
    .S(_05996_),
    .X(_05999_));
 sky130_fd_sc_hd__clkbuf_1 _11980_ (.A(_05999_),
    .X(_00481_));
 sky130_fd_sc_hd__mux2_1 _11981_ (.A0(\regs[5][3] ),
    .A1(_05823_),
    .S(_05996_),
    .X(_06000_));
 sky130_fd_sc_hd__clkbuf_1 _11982_ (.A(_06000_),
    .X(_00482_));
 sky130_fd_sc_hd__mux2_1 _11983_ (.A0(\regs[5][4] ),
    .A1(_05825_),
    .S(_05996_),
    .X(_06001_));
 sky130_fd_sc_hd__clkbuf_1 _11984_ (.A(_06001_),
    .X(_00483_));
 sky130_fd_sc_hd__mux2_1 _11985_ (.A0(\regs[5][5] ),
    .A1(_05827_),
    .S(_05996_),
    .X(_06002_));
 sky130_fd_sc_hd__clkbuf_1 _11986_ (.A(_06002_),
    .X(_00484_));
 sky130_fd_sc_hd__mux2_1 _11987_ (.A0(\regs[5][6] ),
    .A1(_05829_),
    .S(_05996_),
    .X(_06003_));
 sky130_fd_sc_hd__clkbuf_1 _11988_ (.A(_06003_),
    .X(_00485_));
 sky130_fd_sc_hd__mux2_1 _11989_ (.A0(\regs[5][7] ),
    .A1(_05831_),
    .S(_05996_),
    .X(_06004_));
 sky130_fd_sc_hd__clkbuf_1 _11990_ (.A(_06004_),
    .X(_00486_));
 sky130_fd_sc_hd__mux2_1 _11991_ (.A0(\regs[5][8] ),
    .A1(_05833_),
    .S(_05996_),
    .X(_06005_));
 sky130_fd_sc_hd__clkbuf_1 _11992_ (.A(_06005_),
    .X(_00487_));
 sky130_fd_sc_hd__mux2_1 _11993_ (.A0(\regs[5][9] ),
    .A1(_05835_),
    .S(_05996_),
    .X(_06006_));
 sky130_fd_sc_hd__clkbuf_1 _11994_ (.A(_06006_),
    .X(_00488_));
 sky130_fd_sc_hd__clkbuf_8 _11995_ (.A(_05995_),
    .X(_06007_));
 sky130_fd_sc_hd__mux2_1 _11996_ (.A0(\regs[5][10] ),
    .A1(_05837_),
    .S(_06007_),
    .X(_06008_));
 sky130_fd_sc_hd__clkbuf_1 _11997_ (.A(_06008_),
    .X(_00489_));
 sky130_fd_sc_hd__mux2_1 _11998_ (.A0(\regs[5][11] ),
    .A1(_05840_),
    .S(_06007_),
    .X(_06009_));
 sky130_fd_sc_hd__clkbuf_1 _11999_ (.A(_06009_),
    .X(_00490_));
 sky130_fd_sc_hd__mux2_1 _12000_ (.A0(\regs[5][12] ),
    .A1(_05842_),
    .S(_06007_),
    .X(_06010_));
 sky130_fd_sc_hd__clkbuf_1 _12001_ (.A(_06010_),
    .X(_00491_));
 sky130_fd_sc_hd__mux2_1 _12002_ (.A0(\regs[5][13] ),
    .A1(_05844_),
    .S(_06007_),
    .X(_06011_));
 sky130_fd_sc_hd__clkbuf_1 _12003_ (.A(_06011_),
    .X(_00492_));
 sky130_fd_sc_hd__mux2_1 _12004_ (.A0(\regs[5][14] ),
    .A1(_05846_),
    .S(_06007_),
    .X(_06012_));
 sky130_fd_sc_hd__clkbuf_1 _12005_ (.A(_06012_),
    .X(_00493_));
 sky130_fd_sc_hd__mux2_1 _12006_ (.A0(\regs[5][15] ),
    .A1(_05848_),
    .S(_06007_),
    .X(_06013_));
 sky130_fd_sc_hd__clkbuf_1 _12007_ (.A(_06013_),
    .X(_00494_));
 sky130_fd_sc_hd__mux2_1 _12008_ (.A0(\regs[5][16] ),
    .A1(_05850_),
    .S(_06007_),
    .X(_06014_));
 sky130_fd_sc_hd__clkbuf_1 _12009_ (.A(_06014_),
    .X(_00495_));
 sky130_fd_sc_hd__mux2_1 _12010_ (.A0(\regs[5][17] ),
    .A1(_05852_),
    .S(_06007_),
    .X(_06015_));
 sky130_fd_sc_hd__clkbuf_1 _12011_ (.A(_06015_),
    .X(_00496_));
 sky130_fd_sc_hd__mux2_1 _12012_ (.A0(\regs[5][18] ),
    .A1(_05854_),
    .S(_06007_),
    .X(_06016_));
 sky130_fd_sc_hd__clkbuf_1 _12013_ (.A(_06016_),
    .X(_00497_));
 sky130_fd_sc_hd__mux2_1 _12014_ (.A0(\regs[5][19] ),
    .A1(_05856_),
    .S(_06007_),
    .X(_06017_));
 sky130_fd_sc_hd__clkbuf_1 _12015_ (.A(_06017_),
    .X(_00498_));
 sky130_fd_sc_hd__buf_8 _12016_ (.A(_05995_),
    .X(_06018_));
 sky130_fd_sc_hd__mux2_1 _12017_ (.A0(\regs[5][20] ),
    .A1(_05858_),
    .S(_06018_),
    .X(_06019_));
 sky130_fd_sc_hd__clkbuf_1 _12018_ (.A(_06019_),
    .X(_00499_));
 sky130_fd_sc_hd__mux2_1 _12019_ (.A0(\regs[5][21] ),
    .A1(_05861_),
    .S(_06018_),
    .X(_06020_));
 sky130_fd_sc_hd__clkbuf_1 _12020_ (.A(_06020_),
    .X(_00500_));
 sky130_fd_sc_hd__mux2_1 _12021_ (.A0(\regs[5][22] ),
    .A1(_05863_),
    .S(_06018_),
    .X(_06021_));
 sky130_fd_sc_hd__clkbuf_1 _12022_ (.A(_06021_),
    .X(_00501_));
 sky130_fd_sc_hd__mux2_1 _12023_ (.A0(\regs[5][23] ),
    .A1(_05865_),
    .S(_06018_),
    .X(_06022_));
 sky130_fd_sc_hd__clkbuf_1 _12024_ (.A(_06022_),
    .X(_00502_));
 sky130_fd_sc_hd__mux2_1 _12025_ (.A0(\regs[5][24] ),
    .A1(_05867_),
    .S(_06018_),
    .X(_06023_));
 sky130_fd_sc_hd__clkbuf_1 _12026_ (.A(_06023_),
    .X(_00503_));
 sky130_fd_sc_hd__mux2_1 _12027_ (.A0(\regs[5][25] ),
    .A1(_05869_),
    .S(_06018_),
    .X(_06024_));
 sky130_fd_sc_hd__clkbuf_1 _12028_ (.A(_06024_),
    .X(_00504_));
 sky130_fd_sc_hd__mux2_1 _12029_ (.A0(\regs[5][26] ),
    .A1(_05871_),
    .S(_06018_),
    .X(_06025_));
 sky130_fd_sc_hd__clkbuf_1 _12030_ (.A(_06025_),
    .X(_00505_));
 sky130_fd_sc_hd__mux2_1 _12031_ (.A0(\regs[5][27] ),
    .A1(_05873_),
    .S(_06018_),
    .X(_06026_));
 sky130_fd_sc_hd__clkbuf_1 _12032_ (.A(_06026_),
    .X(_00506_));
 sky130_fd_sc_hd__mux2_1 _12033_ (.A0(\regs[5][28] ),
    .A1(_05875_),
    .S(_06018_),
    .X(_06027_));
 sky130_fd_sc_hd__clkbuf_1 _12034_ (.A(_06027_),
    .X(_00507_));
 sky130_fd_sc_hd__mux2_1 _12035_ (.A0(\regs[5][29] ),
    .A1(_05877_),
    .S(_06018_),
    .X(_06028_));
 sky130_fd_sc_hd__clkbuf_1 _12036_ (.A(_06028_),
    .X(_00508_));
 sky130_fd_sc_hd__mux2_1 _12037_ (.A0(\regs[5][30] ),
    .A1(_05879_),
    .S(_05995_),
    .X(_06029_));
 sky130_fd_sc_hd__clkbuf_1 _12038_ (.A(_06029_),
    .X(_00509_));
 sky130_fd_sc_hd__mux2_1 _12039_ (.A0(\regs[5][31] ),
    .A1(_05881_),
    .S(_05995_),
    .X(_06030_));
 sky130_fd_sc_hd__clkbuf_1 _12040_ (.A(_06030_),
    .X(_00510_));
 sky130_fd_sc_hd__o21ai_4 _12041_ (.A1(_01648_),
    .A2(_01642_),
    .B1(_04765_),
    .Y(_06031_));
 sky130_fd_sc_hd__nand2_4 _12042_ (.A(_04767_),
    .B(_06031_),
    .Y(_06032_));
 sky130_fd_sc_hd__buf_6 _12043_ (.A(_06032_),
    .X(_06033_));
 sky130_fd_sc_hd__mux2_1 _12044_ (.A0(_04762_),
    .A1(\regs[8][0] ),
    .S(_06033_),
    .X(_06034_));
 sky130_fd_sc_hd__clkbuf_1 _12045_ (.A(_06034_),
    .X(_00511_));
 sky130_fd_sc_hd__mux2_1 _12046_ (.A0(_04818_),
    .A1(\regs[8][1] ),
    .S(_06033_),
    .X(_06035_));
 sky130_fd_sc_hd__clkbuf_1 _12047_ (.A(_06035_),
    .X(_00512_));
 sky130_fd_sc_hd__mux2_1 _12048_ (.A0(_04858_),
    .A1(\regs[8][2] ),
    .S(_06033_),
    .X(_06036_));
 sky130_fd_sc_hd__clkbuf_1 _12049_ (.A(_06036_),
    .X(_00513_));
 sky130_fd_sc_hd__mux2_1 _12050_ (.A0(_04904_),
    .A1(\regs[8][3] ),
    .S(_06033_),
    .X(_06037_));
 sky130_fd_sc_hd__clkbuf_1 _12051_ (.A(_06037_),
    .X(_00514_));
 sky130_fd_sc_hd__mux2_1 _12052_ (.A0(_04952_),
    .A1(\regs[8][4] ),
    .S(_06033_),
    .X(_06038_));
 sky130_fd_sc_hd__clkbuf_1 _12053_ (.A(_06038_),
    .X(_00515_));
 sky130_fd_sc_hd__mux2_1 _12054_ (.A0(_04992_),
    .A1(\regs[8][5] ),
    .S(_06033_),
    .X(_06039_));
 sky130_fd_sc_hd__clkbuf_1 _12055_ (.A(_06039_),
    .X(_00516_));
 sky130_fd_sc_hd__mux2_1 _12056_ (.A0(_05030_),
    .A1(\regs[8][6] ),
    .S(_06033_),
    .X(_06040_));
 sky130_fd_sc_hd__clkbuf_1 _12057_ (.A(_06040_),
    .X(_00517_));
 sky130_fd_sc_hd__mux2_1 _12058_ (.A0(_05080_),
    .A1(\regs[8][7] ),
    .S(_06033_),
    .X(_06041_));
 sky130_fd_sc_hd__clkbuf_1 _12059_ (.A(_06041_),
    .X(_00518_));
 sky130_fd_sc_hd__mux2_1 _12060_ (.A0(_05121_),
    .A1(\regs[8][8] ),
    .S(_06033_),
    .X(_06042_));
 sky130_fd_sc_hd__clkbuf_1 _12061_ (.A(_06042_),
    .X(_00519_));
 sky130_fd_sc_hd__mux2_1 _12062_ (.A0(_05157_),
    .A1(\regs[8][9] ),
    .S(_06033_),
    .X(_06043_));
 sky130_fd_sc_hd__clkbuf_1 _12063_ (.A(_06043_),
    .X(_00520_));
 sky130_fd_sc_hd__buf_4 _12064_ (.A(_06032_),
    .X(_06044_));
 sky130_fd_sc_hd__mux2_1 _12065_ (.A0(_05187_),
    .A1(\regs[8][10] ),
    .S(_06044_),
    .X(_06045_));
 sky130_fd_sc_hd__clkbuf_1 _12066_ (.A(_06045_),
    .X(_00521_));
 sky130_fd_sc_hd__mux2_1 _12067_ (.A0(_05224_),
    .A1(\regs[8][11] ),
    .S(_06044_),
    .X(_06046_));
 sky130_fd_sc_hd__clkbuf_1 _12068_ (.A(_06046_),
    .X(_00522_));
 sky130_fd_sc_hd__mux2_1 _12069_ (.A0(_05263_),
    .A1(\regs[8][12] ),
    .S(_06044_),
    .X(_06047_));
 sky130_fd_sc_hd__clkbuf_1 _12070_ (.A(_06047_),
    .X(_00523_));
 sky130_fd_sc_hd__mux2_1 _12071_ (.A0(_05296_),
    .A1(\regs[8][13] ),
    .S(_06044_),
    .X(_06048_));
 sky130_fd_sc_hd__clkbuf_1 _12072_ (.A(_06048_),
    .X(_00524_));
 sky130_fd_sc_hd__mux2_1 _12073_ (.A0(_05329_),
    .A1(\regs[8][14] ),
    .S(_06044_),
    .X(_06049_));
 sky130_fd_sc_hd__clkbuf_1 _12074_ (.A(_06049_),
    .X(_00525_));
 sky130_fd_sc_hd__mux2_1 _12075_ (.A0(_05359_),
    .A1(\regs[8][15] ),
    .S(_06044_),
    .X(_06050_));
 sky130_fd_sc_hd__clkbuf_1 _12076_ (.A(_06050_),
    .X(_00526_));
 sky130_fd_sc_hd__mux2_1 _12077_ (.A0(_05400_),
    .A1(\regs[8][16] ),
    .S(_06044_),
    .X(_06051_));
 sky130_fd_sc_hd__clkbuf_1 _12078_ (.A(_06051_),
    .X(_00527_));
 sky130_fd_sc_hd__mux2_1 _12079_ (.A0(_05424_),
    .A1(\regs[8][17] ),
    .S(_06044_),
    .X(_06052_));
 sky130_fd_sc_hd__clkbuf_1 _12080_ (.A(_06052_),
    .X(_00528_));
 sky130_fd_sc_hd__mux2_1 _12081_ (.A0(_05452_),
    .A1(\regs[8][18] ),
    .S(_06044_),
    .X(_06053_));
 sky130_fd_sc_hd__clkbuf_1 _12082_ (.A(_06053_),
    .X(_00529_));
 sky130_fd_sc_hd__mux2_1 _12083_ (.A0(_05477_),
    .A1(\regs[8][19] ),
    .S(_06044_),
    .X(_06054_));
 sky130_fd_sc_hd__clkbuf_1 _12084_ (.A(_06054_),
    .X(_00530_));
 sky130_fd_sc_hd__buf_8 _12085_ (.A(_06032_),
    .X(_06055_));
 sky130_fd_sc_hd__mux2_1 _12086_ (.A0(_05514_),
    .A1(\regs[8][20] ),
    .S(_06055_),
    .X(_06056_));
 sky130_fd_sc_hd__clkbuf_1 _12087_ (.A(_06056_),
    .X(_00531_));
 sky130_fd_sc_hd__mux2_1 _12088_ (.A0(_05541_),
    .A1(\regs[8][21] ),
    .S(_06055_),
    .X(_06057_));
 sky130_fd_sc_hd__clkbuf_1 _12089_ (.A(_06057_),
    .X(_00532_));
 sky130_fd_sc_hd__mux2_1 _12090_ (.A0(_05570_),
    .A1(\regs[8][22] ),
    .S(_06055_),
    .X(_06058_));
 sky130_fd_sc_hd__clkbuf_1 _12091_ (.A(_06058_),
    .X(_00533_));
 sky130_fd_sc_hd__mux2_1 _12092_ (.A0(_05600_),
    .A1(\regs[8][23] ),
    .S(_06055_),
    .X(_06059_));
 sky130_fd_sc_hd__clkbuf_1 _12093_ (.A(_06059_),
    .X(_00534_));
 sky130_fd_sc_hd__mux2_1 _12094_ (.A0(_05636_),
    .A1(\regs[8][24] ),
    .S(_06055_),
    .X(_06060_));
 sky130_fd_sc_hd__clkbuf_1 _12095_ (.A(_06060_),
    .X(_00535_));
 sky130_fd_sc_hd__mux2_1 _12096_ (.A0(_05660_),
    .A1(\regs[8][25] ),
    .S(_06055_),
    .X(_06061_));
 sky130_fd_sc_hd__clkbuf_1 _12097_ (.A(_06061_),
    .X(_00536_));
 sky130_fd_sc_hd__mux2_1 _12098_ (.A0(_05684_),
    .A1(\regs[8][26] ),
    .S(_06055_),
    .X(_06062_));
 sky130_fd_sc_hd__clkbuf_1 _12099_ (.A(_06062_),
    .X(_00537_));
 sky130_fd_sc_hd__mux2_1 _12100_ (.A0(_05708_),
    .A1(\regs[8][27] ),
    .S(_06055_),
    .X(_06063_));
 sky130_fd_sc_hd__clkbuf_1 _12101_ (.A(_06063_),
    .X(_00538_));
 sky130_fd_sc_hd__mux2_1 _12102_ (.A0(_05735_),
    .A1(\regs[8][28] ),
    .S(_06055_),
    .X(_06064_));
 sky130_fd_sc_hd__clkbuf_1 _12103_ (.A(_06064_),
    .X(_00539_));
 sky130_fd_sc_hd__mux2_1 _12104_ (.A0(_05763_),
    .A1(\regs[8][29] ),
    .S(_06055_),
    .X(_06065_));
 sky130_fd_sc_hd__clkbuf_1 _12105_ (.A(_06065_),
    .X(_00540_));
 sky130_fd_sc_hd__mux2_1 _12106_ (.A0(_05787_),
    .A1(\regs[8][30] ),
    .S(_06032_),
    .X(_06066_));
 sky130_fd_sc_hd__clkbuf_1 _12107_ (.A(_06066_),
    .X(_00541_));
 sky130_fd_sc_hd__mux2_1 _12108_ (.A0(_05811_),
    .A1(\regs[8][31] ),
    .S(_06032_),
    .X(_06067_));
 sky130_fd_sc_hd__clkbuf_1 _12109_ (.A(_06067_),
    .X(_00542_));
 sky130_fd_sc_hd__clkinv_2 _12110_ (.A(_04755_),
    .Y(_06068_));
 sky130_fd_sc_hd__buf_6 _12111_ (.A(_06068_),
    .X(_00068_));
 sky130_fd_sc_hd__buf_6 _12112_ (.A(_04755_),
    .X(_06069_));
 sky130_fd_sc_hd__buf_6 _12113_ (.A(_06069_),
    .X(_06070_));
 sky130_fd_sc_hd__inv_2 _12114_ (.A(_06070_),
    .Y(_00069_));
 sky130_fd_sc_hd__inv_2 _12115_ (.A(_06070_),
    .Y(_00070_));
 sky130_fd_sc_hd__inv_2 _12116_ (.A(_06070_),
    .Y(_00071_));
 sky130_fd_sc_hd__or2_1 _12117_ (.A(_01648_),
    .B(_04763_),
    .X(_06071_));
 sky130_fd_sc_hd__clkbuf_4 _12118_ (.A(_06071_),
    .X(_06072_));
 sky130_fd_sc_hd__nor2_4 _12119_ (.A(_06072_),
    .B(_05921_),
    .Y(_06073_));
 sky130_fd_sc_hd__clkbuf_8 _12120_ (.A(_06073_),
    .X(_06074_));
 sky130_fd_sc_hd__mux2_1 _12121_ (.A0(\regs[13][0] ),
    .A1(_05813_),
    .S(_06074_),
    .X(_06075_));
 sky130_fd_sc_hd__clkbuf_1 _12122_ (.A(_06075_),
    .X(_00543_));
 sky130_fd_sc_hd__mux2_1 _12123_ (.A0(\regs[13][1] ),
    .A1(_05819_),
    .S(_06074_),
    .X(_06076_));
 sky130_fd_sc_hd__clkbuf_1 _12124_ (.A(_06076_),
    .X(_00544_));
 sky130_fd_sc_hd__mux2_1 _12125_ (.A0(\regs[13][2] ),
    .A1(_05821_),
    .S(_06074_),
    .X(_06077_));
 sky130_fd_sc_hd__clkbuf_1 _12126_ (.A(_06077_),
    .X(_00545_));
 sky130_fd_sc_hd__mux2_1 _12127_ (.A0(\regs[13][3] ),
    .A1(_05823_),
    .S(_06074_),
    .X(_06078_));
 sky130_fd_sc_hd__clkbuf_1 _12128_ (.A(_06078_),
    .X(_00546_));
 sky130_fd_sc_hd__mux2_1 _12129_ (.A0(\regs[13][4] ),
    .A1(_05825_),
    .S(_06074_),
    .X(_06079_));
 sky130_fd_sc_hd__clkbuf_1 _12130_ (.A(_06079_),
    .X(_00547_));
 sky130_fd_sc_hd__mux2_1 _12131_ (.A0(\regs[13][5] ),
    .A1(_05827_),
    .S(_06074_),
    .X(_06080_));
 sky130_fd_sc_hd__clkbuf_1 _12132_ (.A(_06080_),
    .X(_00548_));
 sky130_fd_sc_hd__mux2_1 _12133_ (.A0(\regs[13][6] ),
    .A1(_05829_),
    .S(_06074_),
    .X(_06081_));
 sky130_fd_sc_hd__clkbuf_1 _12134_ (.A(_06081_),
    .X(_00549_));
 sky130_fd_sc_hd__mux2_1 _12135_ (.A0(\regs[13][7] ),
    .A1(_05831_),
    .S(_06074_),
    .X(_06082_));
 sky130_fd_sc_hd__clkbuf_1 _12136_ (.A(_06082_),
    .X(_00550_));
 sky130_fd_sc_hd__mux2_1 _12137_ (.A0(\regs[13][8] ),
    .A1(_05833_),
    .S(_06074_),
    .X(_06083_));
 sky130_fd_sc_hd__clkbuf_1 _12138_ (.A(_06083_),
    .X(_00551_));
 sky130_fd_sc_hd__mux2_1 _12139_ (.A0(\regs[13][9] ),
    .A1(_05835_),
    .S(_06074_),
    .X(_06084_));
 sky130_fd_sc_hd__clkbuf_1 _12140_ (.A(_06084_),
    .X(_00552_));
 sky130_fd_sc_hd__buf_4 _12141_ (.A(_06073_),
    .X(_06085_));
 sky130_fd_sc_hd__mux2_1 _12142_ (.A0(\regs[13][10] ),
    .A1(_05837_),
    .S(_06085_),
    .X(_06086_));
 sky130_fd_sc_hd__clkbuf_1 _12143_ (.A(_06086_),
    .X(_00553_));
 sky130_fd_sc_hd__mux2_1 _12144_ (.A0(\regs[13][11] ),
    .A1(_05840_),
    .S(_06085_),
    .X(_06087_));
 sky130_fd_sc_hd__clkbuf_1 _12145_ (.A(_06087_),
    .X(_00554_));
 sky130_fd_sc_hd__mux2_1 _12146_ (.A0(\regs[13][12] ),
    .A1(_05842_),
    .S(_06085_),
    .X(_06088_));
 sky130_fd_sc_hd__clkbuf_1 _12147_ (.A(_06088_),
    .X(_00555_));
 sky130_fd_sc_hd__mux2_1 _12148_ (.A0(\regs[13][13] ),
    .A1(_05844_),
    .S(_06085_),
    .X(_06089_));
 sky130_fd_sc_hd__clkbuf_1 _12149_ (.A(_06089_),
    .X(_00556_));
 sky130_fd_sc_hd__mux2_1 _12150_ (.A0(\regs[13][14] ),
    .A1(_05846_),
    .S(_06085_),
    .X(_06090_));
 sky130_fd_sc_hd__clkbuf_1 _12151_ (.A(_06090_),
    .X(_00557_));
 sky130_fd_sc_hd__mux2_1 _12152_ (.A0(\regs[13][15] ),
    .A1(_05848_),
    .S(_06085_),
    .X(_06091_));
 sky130_fd_sc_hd__clkbuf_1 _12153_ (.A(_06091_),
    .X(_00558_));
 sky130_fd_sc_hd__mux2_1 _12154_ (.A0(\regs[13][16] ),
    .A1(_05850_),
    .S(_06085_),
    .X(_06092_));
 sky130_fd_sc_hd__clkbuf_1 _12155_ (.A(_06092_),
    .X(_00559_));
 sky130_fd_sc_hd__mux2_1 _12156_ (.A0(\regs[13][17] ),
    .A1(_05852_),
    .S(_06085_),
    .X(_06093_));
 sky130_fd_sc_hd__clkbuf_1 _12157_ (.A(_06093_),
    .X(_00560_));
 sky130_fd_sc_hd__mux2_1 _12158_ (.A0(\regs[13][18] ),
    .A1(_05854_),
    .S(_06085_),
    .X(_06094_));
 sky130_fd_sc_hd__clkbuf_1 _12159_ (.A(_06094_),
    .X(_00561_));
 sky130_fd_sc_hd__mux2_1 _12160_ (.A0(\regs[13][19] ),
    .A1(_05856_),
    .S(_06085_),
    .X(_06095_));
 sky130_fd_sc_hd__clkbuf_1 _12161_ (.A(_06095_),
    .X(_00562_));
 sky130_fd_sc_hd__buf_6 _12162_ (.A(_06073_),
    .X(_06096_));
 sky130_fd_sc_hd__mux2_1 _12163_ (.A0(\regs[13][20] ),
    .A1(_05858_),
    .S(_06096_),
    .X(_06097_));
 sky130_fd_sc_hd__clkbuf_1 _12164_ (.A(_06097_),
    .X(_00563_));
 sky130_fd_sc_hd__mux2_1 _12165_ (.A0(\regs[13][21] ),
    .A1(_05861_),
    .S(_06096_),
    .X(_06098_));
 sky130_fd_sc_hd__clkbuf_1 _12166_ (.A(_06098_),
    .X(_00564_));
 sky130_fd_sc_hd__mux2_1 _12167_ (.A0(\regs[13][22] ),
    .A1(_05863_),
    .S(_06096_),
    .X(_06099_));
 sky130_fd_sc_hd__clkbuf_1 _12168_ (.A(_06099_),
    .X(_00565_));
 sky130_fd_sc_hd__mux2_1 _12169_ (.A0(\regs[13][23] ),
    .A1(_05865_),
    .S(_06096_),
    .X(_06100_));
 sky130_fd_sc_hd__clkbuf_1 _12170_ (.A(_06100_),
    .X(_00566_));
 sky130_fd_sc_hd__mux2_1 _12171_ (.A0(\regs[13][24] ),
    .A1(_05867_),
    .S(_06096_),
    .X(_06101_));
 sky130_fd_sc_hd__clkbuf_1 _12172_ (.A(_06101_),
    .X(_00567_));
 sky130_fd_sc_hd__mux2_1 _12173_ (.A0(\regs[13][25] ),
    .A1(_05869_),
    .S(_06096_),
    .X(_06102_));
 sky130_fd_sc_hd__clkbuf_1 _12174_ (.A(_06102_),
    .X(_00568_));
 sky130_fd_sc_hd__mux2_1 _12175_ (.A0(\regs[13][26] ),
    .A1(_05871_),
    .S(_06096_),
    .X(_06103_));
 sky130_fd_sc_hd__clkbuf_1 _12176_ (.A(_06103_),
    .X(_00569_));
 sky130_fd_sc_hd__mux2_1 _12177_ (.A0(\regs[13][27] ),
    .A1(_05873_),
    .S(_06096_),
    .X(_06104_));
 sky130_fd_sc_hd__clkbuf_1 _12178_ (.A(_06104_),
    .X(_00570_));
 sky130_fd_sc_hd__mux2_1 _12179_ (.A0(\regs[13][28] ),
    .A1(_05875_),
    .S(_06096_),
    .X(_06105_));
 sky130_fd_sc_hd__clkbuf_1 _12180_ (.A(_06105_),
    .X(_00571_));
 sky130_fd_sc_hd__mux2_1 _12181_ (.A0(\regs[13][29] ),
    .A1(_05877_),
    .S(_06096_),
    .X(_06106_));
 sky130_fd_sc_hd__clkbuf_1 _12182_ (.A(_06106_),
    .X(_00572_));
 sky130_fd_sc_hd__mux2_1 _12183_ (.A0(\regs[13][30] ),
    .A1(_05879_),
    .S(_06073_),
    .X(_06107_));
 sky130_fd_sc_hd__clkbuf_1 _12184_ (.A(_06107_),
    .X(_00573_));
 sky130_fd_sc_hd__mux2_1 _12185_ (.A0(\regs[13][31] ),
    .A1(_05881_),
    .S(_06073_),
    .X(_06108_));
 sky130_fd_sc_hd__clkbuf_1 _12186_ (.A(_06108_),
    .X(_00574_));
 sky130_fd_sc_hd__nor2_4 _12187_ (.A(_05883_),
    .B(_05921_),
    .Y(_06109_));
 sky130_fd_sc_hd__clkbuf_8 _12188_ (.A(_06109_),
    .X(_06110_));
 sky130_fd_sc_hd__mux2_1 _12189_ (.A0(\regs[14][0] ),
    .A1(_05813_),
    .S(_06110_),
    .X(_06111_));
 sky130_fd_sc_hd__clkbuf_1 _12190_ (.A(_06111_),
    .X(_00575_));
 sky130_fd_sc_hd__mux2_1 _12191_ (.A0(\regs[14][1] ),
    .A1(_05819_),
    .S(_06110_),
    .X(_06112_));
 sky130_fd_sc_hd__clkbuf_1 _12192_ (.A(_06112_),
    .X(_00576_));
 sky130_fd_sc_hd__mux2_1 _12193_ (.A0(\regs[14][2] ),
    .A1(_05821_),
    .S(_06110_),
    .X(_06113_));
 sky130_fd_sc_hd__clkbuf_1 _12194_ (.A(_06113_),
    .X(_00577_));
 sky130_fd_sc_hd__mux2_1 _12195_ (.A0(\regs[14][3] ),
    .A1(_05823_),
    .S(_06110_),
    .X(_06114_));
 sky130_fd_sc_hd__clkbuf_1 _12196_ (.A(_06114_),
    .X(_00578_));
 sky130_fd_sc_hd__mux2_1 _12197_ (.A0(\regs[14][4] ),
    .A1(_05825_),
    .S(_06110_),
    .X(_06115_));
 sky130_fd_sc_hd__clkbuf_1 _12198_ (.A(_06115_),
    .X(_00579_));
 sky130_fd_sc_hd__mux2_1 _12199_ (.A0(\regs[14][5] ),
    .A1(_05827_),
    .S(_06110_),
    .X(_06116_));
 sky130_fd_sc_hd__clkbuf_1 _12200_ (.A(_06116_),
    .X(_00580_));
 sky130_fd_sc_hd__mux2_1 _12201_ (.A0(\regs[14][6] ),
    .A1(_05829_),
    .S(_06110_),
    .X(_06117_));
 sky130_fd_sc_hd__clkbuf_1 _12202_ (.A(_06117_),
    .X(_00581_));
 sky130_fd_sc_hd__mux2_1 _12203_ (.A0(\regs[14][7] ),
    .A1(_05831_),
    .S(_06110_),
    .X(_06118_));
 sky130_fd_sc_hd__clkbuf_1 _12204_ (.A(_06118_),
    .X(_00582_));
 sky130_fd_sc_hd__mux2_1 _12205_ (.A0(\regs[14][8] ),
    .A1(_05833_),
    .S(_06110_),
    .X(_06119_));
 sky130_fd_sc_hd__clkbuf_1 _12206_ (.A(_06119_),
    .X(_00583_));
 sky130_fd_sc_hd__mux2_1 _12207_ (.A0(\regs[14][9] ),
    .A1(_05835_),
    .S(_06110_),
    .X(_06120_));
 sky130_fd_sc_hd__clkbuf_1 _12208_ (.A(_06120_),
    .X(_00584_));
 sky130_fd_sc_hd__buf_4 _12209_ (.A(_06109_),
    .X(_06121_));
 sky130_fd_sc_hd__mux2_1 _12210_ (.A0(\regs[14][10] ),
    .A1(_05837_),
    .S(_06121_),
    .X(_06122_));
 sky130_fd_sc_hd__clkbuf_1 _12211_ (.A(_06122_),
    .X(_00585_));
 sky130_fd_sc_hd__mux2_1 _12212_ (.A0(\regs[14][11] ),
    .A1(_05840_),
    .S(_06121_),
    .X(_06123_));
 sky130_fd_sc_hd__clkbuf_1 _12213_ (.A(_06123_),
    .X(_00586_));
 sky130_fd_sc_hd__mux2_1 _12214_ (.A0(\regs[14][12] ),
    .A1(_05842_),
    .S(_06121_),
    .X(_06124_));
 sky130_fd_sc_hd__clkbuf_1 _12215_ (.A(_06124_),
    .X(_00587_));
 sky130_fd_sc_hd__mux2_1 _12216_ (.A0(\regs[14][13] ),
    .A1(_05844_),
    .S(_06121_),
    .X(_06125_));
 sky130_fd_sc_hd__clkbuf_1 _12217_ (.A(_06125_),
    .X(_00588_));
 sky130_fd_sc_hd__mux2_1 _12218_ (.A0(\regs[14][14] ),
    .A1(_05846_),
    .S(_06121_),
    .X(_06126_));
 sky130_fd_sc_hd__clkbuf_1 _12219_ (.A(_06126_),
    .X(_00589_));
 sky130_fd_sc_hd__mux2_1 _12220_ (.A0(\regs[14][15] ),
    .A1(_05848_),
    .S(_06121_),
    .X(_06127_));
 sky130_fd_sc_hd__clkbuf_1 _12221_ (.A(_06127_),
    .X(_00590_));
 sky130_fd_sc_hd__mux2_1 _12222_ (.A0(\regs[14][16] ),
    .A1(_05850_),
    .S(_06121_),
    .X(_06128_));
 sky130_fd_sc_hd__clkbuf_1 _12223_ (.A(_06128_),
    .X(_00591_));
 sky130_fd_sc_hd__mux2_1 _12224_ (.A0(\regs[14][17] ),
    .A1(_05852_),
    .S(_06121_),
    .X(_06129_));
 sky130_fd_sc_hd__clkbuf_1 _12225_ (.A(_06129_),
    .X(_00592_));
 sky130_fd_sc_hd__mux2_1 _12226_ (.A0(\regs[14][18] ),
    .A1(_05854_),
    .S(_06121_),
    .X(_06130_));
 sky130_fd_sc_hd__clkbuf_1 _12227_ (.A(_06130_),
    .X(_00593_));
 sky130_fd_sc_hd__mux2_1 _12228_ (.A0(\regs[14][19] ),
    .A1(_05856_),
    .S(_06121_),
    .X(_06131_));
 sky130_fd_sc_hd__clkbuf_1 _12229_ (.A(_06131_),
    .X(_00594_));
 sky130_fd_sc_hd__buf_6 _12230_ (.A(_06109_),
    .X(_06132_));
 sky130_fd_sc_hd__mux2_1 _12231_ (.A0(\regs[14][20] ),
    .A1(_05858_),
    .S(_06132_),
    .X(_06133_));
 sky130_fd_sc_hd__clkbuf_1 _12232_ (.A(_06133_),
    .X(_00595_));
 sky130_fd_sc_hd__mux2_1 _12233_ (.A0(\regs[14][21] ),
    .A1(_05861_),
    .S(_06132_),
    .X(_06134_));
 sky130_fd_sc_hd__clkbuf_1 _12234_ (.A(_06134_),
    .X(_00596_));
 sky130_fd_sc_hd__mux2_1 _12235_ (.A0(\regs[14][22] ),
    .A1(_05863_),
    .S(_06132_),
    .X(_06135_));
 sky130_fd_sc_hd__clkbuf_1 _12236_ (.A(_06135_),
    .X(_00597_));
 sky130_fd_sc_hd__mux2_1 _12237_ (.A0(\regs[14][23] ),
    .A1(_05865_),
    .S(_06132_),
    .X(_06136_));
 sky130_fd_sc_hd__clkbuf_1 _12238_ (.A(_06136_),
    .X(_00598_));
 sky130_fd_sc_hd__mux2_1 _12239_ (.A0(\regs[14][24] ),
    .A1(_05867_),
    .S(_06132_),
    .X(_06137_));
 sky130_fd_sc_hd__clkbuf_1 _12240_ (.A(_06137_),
    .X(_00599_));
 sky130_fd_sc_hd__mux2_1 _12241_ (.A0(\regs[14][25] ),
    .A1(_05869_),
    .S(_06132_),
    .X(_06138_));
 sky130_fd_sc_hd__clkbuf_1 _12242_ (.A(_06138_),
    .X(_00600_));
 sky130_fd_sc_hd__mux2_1 _12243_ (.A0(\regs[14][26] ),
    .A1(_05871_),
    .S(_06132_),
    .X(_06139_));
 sky130_fd_sc_hd__clkbuf_1 _12244_ (.A(_06139_),
    .X(_00601_));
 sky130_fd_sc_hd__mux2_1 _12245_ (.A0(\regs[14][27] ),
    .A1(_05873_),
    .S(_06132_),
    .X(_06140_));
 sky130_fd_sc_hd__clkbuf_1 _12246_ (.A(_06140_),
    .X(_00602_));
 sky130_fd_sc_hd__mux2_1 _12247_ (.A0(\regs[14][28] ),
    .A1(_05875_),
    .S(_06132_),
    .X(_06141_));
 sky130_fd_sc_hd__clkbuf_1 _12248_ (.A(_06141_),
    .X(_00603_));
 sky130_fd_sc_hd__mux2_1 _12249_ (.A0(\regs[14][29] ),
    .A1(_05877_),
    .S(_06132_),
    .X(_06142_));
 sky130_fd_sc_hd__clkbuf_1 _12250_ (.A(_06142_),
    .X(_00604_));
 sky130_fd_sc_hd__mux2_1 _12251_ (.A0(\regs[14][30] ),
    .A1(_05879_),
    .S(_06109_),
    .X(_06143_));
 sky130_fd_sc_hd__clkbuf_1 _12252_ (.A(_06143_),
    .X(_00605_));
 sky130_fd_sc_hd__mux2_1 _12253_ (.A0(\regs[14][31] ),
    .A1(_05881_),
    .S(_06109_),
    .X(_06144_));
 sky130_fd_sc_hd__clkbuf_1 _12254_ (.A(_06144_),
    .X(_00606_));
 sky130_fd_sc_hd__or4bb_4 _12255_ (.A(_02315_),
    .B(_02241_),
    .C_N(_04765_),
    .D_N(_02313_),
    .X(_06145_));
 sky130_fd_sc_hd__nor2_4 _12256_ (.A(_04758_),
    .B(_06145_),
    .Y(_06146_));
 sky130_fd_sc_hd__buf_6 _12257_ (.A(_06146_),
    .X(_06147_));
 sky130_fd_sc_hd__mux2_1 _12258_ (.A0(\regs[16][0] ),
    .A1(_05813_),
    .S(_06147_),
    .X(_06148_));
 sky130_fd_sc_hd__clkbuf_1 _12259_ (.A(_06148_),
    .X(_00607_));
 sky130_fd_sc_hd__mux2_1 _12260_ (.A0(\regs[16][1] ),
    .A1(_05819_),
    .S(_06147_),
    .X(_06149_));
 sky130_fd_sc_hd__clkbuf_1 _12261_ (.A(_06149_),
    .X(_00608_));
 sky130_fd_sc_hd__mux2_1 _12262_ (.A0(\regs[16][2] ),
    .A1(_05821_),
    .S(_06147_),
    .X(_06150_));
 sky130_fd_sc_hd__clkbuf_1 _12263_ (.A(_06150_),
    .X(_00609_));
 sky130_fd_sc_hd__mux2_1 _12264_ (.A0(\regs[16][3] ),
    .A1(_05823_),
    .S(_06147_),
    .X(_06151_));
 sky130_fd_sc_hd__clkbuf_1 _12265_ (.A(_06151_),
    .X(_00610_));
 sky130_fd_sc_hd__mux2_1 _12266_ (.A0(\regs[16][4] ),
    .A1(_05825_),
    .S(_06147_),
    .X(_06152_));
 sky130_fd_sc_hd__clkbuf_1 _12267_ (.A(_06152_),
    .X(_00611_));
 sky130_fd_sc_hd__mux2_1 _12268_ (.A0(\regs[16][5] ),
    .A1(_05827_),
    .S(_06147_),
    .X(_06153_));
 sky130_fd_sc_hd__clkbuf_1 _12269_ (.A(_06153_),
    .X(_00612_));
 sky130_fd_sc_hd__mux2_1 _12270_ (.A0(\regs[16][6] ),
    .A1(_05829_),
    .S(_06147_),
    .X(_06154_));
 sky130_fd_sc_hd__clkbuf_1 _12271_ (.A(_06154_),
    .X(_00613_));
 sky130_fd_sc_hd__mux2_1 _12272_ (.A0(\regs[16][7] ),
    .A1(_05831_),
    .S(_06147_),
    .X(_06155_));
 sky130_fd_sc_hd__clkbuf_1 _12273_ (.A(_06155_),
    .X(_00614_));
 sky130_fd_sc_hd__mux2_1 _12274_ (.A0(\regs[16][8] ),
    .A1(_05833_),
    .S(_06147_),
    .X(_06156_));
 sky130_fd_sc_hd__clkbuf_1 _12275_ (.A(_06156_),
    .X(_00615_));
 sky130_fd_sc_hd__mux2_1 _12276_ (.A0(\regs[16][9] ),
    .A1(_05835_),
    .S(_06147_),
    .X(_06157_));
 sky130_fd_sc_hd__clkbuf_1 _12277_ (.A(_06157_),
    .X(_00616_));
 sky130_fd_sc_hd__buf_6 _12278_ (.A(_06146_),
    .X(_06158_));
 sky130_fd_sc_hd__mux2_1 _12279_ (.A0(\regs[16][10] ),
    .A1(_05837_),
    .S(_06158_),
    .X(_06159_));
 sky130_fd_sc_hd__clkbuf_1 _12280_ (.A(_06159_),
    .X(_00617_));
 sky130_fd_sc_hd__mux2_1 _12281_ (.A0(\regs[16][11] ),
    .A1(_05840_),
    .S(_06158_),
    .X(_06160_));
 sky130_fd_sc_hd__clkbuf_1 _12282_ (.A(_06160_),
    .X(_00618_));
 sky130_fd_sc_hd__mux2_1 _12283_ (.A0(\regs[16][12] ),
    .A1(_05842_),
    .S(_06158_),
    .X(_06161_));
 sky130_fd_sc_hd__clkbuf_1 _12284_ (.A(_06161_),
    .X(_00619_));
 sky130_fd_sc_hd__mux2_1 _12285_ (.A0(\regs[16][13] ),
    .A1(_05844_),
    .S(_06158_),
    .X(_06162_));
 sky130_fd_sc_hd__clkbuf_1 _12286_ (.A(_06162_),
    .X(_00620_));
 sky130_fd_sc_hd__mux2_1 _12287_ (.A0(\regs[16][14] ),
    .A1(_05846_),
    .S(_06158_),
    .X(_06163_));
 sky130_fd_sc_hd__clkbuf_1 _12288_ (.A(_06163_),
    .X(_00621_));
 sky130_fd_sc_hd__mux2_1 _12289_ (.A0(\regs[16][15] ),
    .A1(_05848_),
    .S(_06158_),
    .X(_06164_));
 sky130_fd_sc_hd__clkbuf_1 _12290_ (.A(_06164_),
    .X(_00622_));
 sky130_fd_sc_hd__mux2_1 _12291_ (.A0(\regs[16][16] ),
    .A1(_05850_),
    .S(_06158_),
    .X(_06165_));
 sky130_fd_sc_hd__clkbuf_1 _12292_ (.A(_06165_),
    .X(_00623_));
 sky130_fd_sc_hd__mux2_1 _12293_ (.A0(\regs[16][17] ),
    .A1(_05852_),
    .S(_06158_),
    .X(_06166_));
 sky130_fd_sc_hd__clkbuf_1 _12294_ (.A(_06166_),
    .X(_00624_));
 sky130_fd_sc_hd__mux2_1 _12295_ (.A0(\regs[16][18] ),
    .A1(_05854_),
    .S(_06158_),
    .X(_06167_));
 sky130_fd_sc_hd__clkbuf_1 _12296_ (.A(_06167_),
    .X(_00625_));
 sky130_fd_sc_hd__mux2_1 _12297_ (.A0(\regs[16][19] ),
    .A1(_05856_),
    .S(_06158_),
    .X(_06168_));
 sky130_fd_sc_hd__clkbuf_1 _12298_ (.A(_06168_),
    .X(_00626_));
 sky130_fd_sc_hd__buf_6 _12299_ (.A(_06146_),
    .X(_06169_));
 sky130_fd_sc_hd__mux2_1 _12300_ (.A0(\regs[16][20] ),
    .A1(_05858_),
    .S(_06169_),
    .X(_06170_));
 sky130_fd_sc_hd__clkbuf_1 _12301_ (.A(_06170_),
    .X(_00627_));
 sky130_fd_sc_hd__mux2_1 _12302_ (.A0(\regs[16][21] ),
    .A1(_05861_),
    .S(_06169_),
    .X(_06171_));
 sky130_fd_sc_hd__clkbuf_1 _12303_ (.A(_06171_),
    .X(_00628_));
 sky130_fd_sc_hd__mux2_1 _12304_ (.A0(\regs[16][22] ),
    .A1(_05863_),
    .S(_06169_),
    .X(_06172_));
 sky130_fd_sc_hd__clkbuf_1 _12305_ (.A(_06172_),
    .X(_00629_));
 sky130_fd_sc_hd__mux2_1 _12306_ (.A0(\regs[16][23] ),
    .A1(_05865_),
    .S(_06169_),
    .X(_06173_));
 sky130_fd_sc_hd__clkbuf_1 _12307_ (.A(_06173_),
    .X(_00630_));
 sky130_fd_sc_hd__mux2_1 _12308_ (.A0(\regs[16][24] ),
    .A1(_05867_),
    .S(_06169_),
    .X(_06174_));
 sky130_fd_sc_hd__clkbuf_1 _12309_ (.A(_06174_),
    .X(_00631_));
 sky130_fd_sc_hd__mux2_1 _12310_ (.A0(\regs[16][25] ),
    .A1(_05869_),
    .S(_06169_),
    .X(_06175_));
 sky130_fd_sc_hd__clkbuf_1 _12311_ (.A(_06175_),
    .X(_00632_));
 sky130_fd_sc_hd__mux2_1 _12312_ (.A0(\regs[16][26] ),
    .A1(_05871_),
    .S(_06169_),
    .X(_06176_));
 sky130_fd_sc_hd__clkbuf_1 _12313_ (.A(_06176_),
    .X(_00633_));
 sky130_fd_sc_hd__mux2_1 _12314_ (.A0(\regs[16][27] ),
    .A1(_05873_),
    .S(_06169_),
    .X(_06177_));
 sky130_fd_sc_hd__clkbuf_1 _12315_ (.A(_06177_),
    .X(_00634_));
 sky130_fd_sc_hd__mux2_1 _12316_ (.A0(\regs[16][28] ),
    .A1(_05875_),
    .S(_06169_),
    .X(_06178_));
 sky130_fd_sc_hd__clkbuf_1 _12317_ (.A(_06178_),
    .X(_00635_));
 sky130_fd_sc_hd__mux2_1 _12318_ (.A0(\regs[16][29] ),
    .A1(_05877_),
    .S(_06169_),
    .X(_06179_));
 sky130_fd_sc_hd__clkbuf_1 _12319_ (.A(_06179_),
    .X(_00636_));
 sky130_fd_sc_hd__mux2_1 _12320_ (.A0(\regs[16][30] ),
    .A1(_05879_),
    .S(_06146_),
    .X(_06180_));
 sky130_fd_sc_hd__clkbuf_1 _12321_ (.A(_06180_),
    .X(_00637_));
 sky130_fd_sc_hd__mux2_1 _12322_ (.A0(\regs[16][31] ),
    .A1(_05881_),
    .S(_06146_),
    .X(_06181_));
 sky130_fd_sc_hd__clkbuf_1 _12323_ (.A(_06181_),
    .X(_00638_));
 sky130_fd_sc_hd__nand2_4 _12324_ (.A(_04767_),
    .B(_05814_),
    .Y(_06182_));
 sky130_fd_sc_hd__clkbuf_8 _12325_ (.A(_06182_),
    .X(_06183_));
 sky130_fd_sc_hd__mux2_1 _12326_ (.A0(_04762_),
    .A1(\regs[11][0] ),
    .S(_06183_),
    .X(_06184_));
 sky130_fd_sc_hd__clkbuf_1 _12327_ (.A(_06184_),
    .X(_00639_));
 sky130_fd_sc_hd__mux2_1 _12328_ (.A0(_04818_),
    .A1(\regs[11][1] ),
    .S(_06183_),
    .X(_06185_));
 sky130_fd_sc_hd__clkbuf_1 _12329_ (.A(_06185_),
    .X(_00640_));
 sky130_fd_sc_hd__mux2_1 _12330_ (.A0(_04858_),
    .A1(\regs[11][2] ),
    .S(_06183_),
    .X(_06186_));
 sky130_fd_sc_hd__clkbuf_1 _12331_ (.A(_06186_),
    .X(_00641_));
 sky130_fd_sc_hd__mux2_1 _12332_ (.A0(_04904_),
    .A1(\regs[11][3] ),
    .S(_06183_),
    .X(_06187_));
 sky130_fd_sc_hd__clkbuf_1 _12333_ (.A(_06187_),
    .X(_00642_));
 sky130_fd_sc_hd__mux2_1 _12334_ (.A0(_04952_),
    .A1(\regs[11][4] ),
    .S(_06183_),
    .X(_06188_));
 sky130_fd_sc_hd__clkbuf_1 _12335_ (.A(_06188_),
    .X(_00643_));
 sky130_fd_sc_hd__mux2_1 _12336_ (.A0(_04992_),
    .A1(\regs[11][5] ),
    .S(_06183_),
    .X(_06189_));
 sky130_fd_sc_hd__clkbuf_1 _12337_ (.A(_06189_),
    .X(_00644_));
 sky130_fd_sc_hd__mux2_1 _12338_ (.A0(_05030_),
    .A1(\regs[11][6] ),
    .S(_06183_),
    .X(_06190_));
 sky130_fd_sc_hd__clkbuf_1 _12339_ (.A(_06190_),
    .X(_00645_));
 sky130_fd_sc_hd__mux2_1 _12340_ (.A0(_05080_),
    .A1(\regs[11][7] ),
    .S(_06183_),
    .X(_06191_));
 sky130_fd_sc_hd__clkbuf_1 _12341_ (.A(_06191_),
    .X(_00646_));
 sky130_fd_sc_hd__mux2_1 _12342_ (.A0(_05121_),
    .A1(\regs[11][8] ),
    .S(_06183_),
    .X(_06192_));
 sky130_fd_sc_hd__clkbuf_1 _12343_ (.A(_06192_),
    .X(_00647_));
 sky130_fd_sc_hd__mux2_1 _12344_ (.A0(_05157_),
    .A1(\regs[11][9] ),
    .S(_06183_),
    .X(_06193_));
 sky130_fd_sc_hd__clkbuf_1 _12345_ (.A(_06193_),
    .X(_00648_));
 sky130_fd_sc_hd__buf_4 _12346_ (.A(_06182_),
    .X(_06194_));
 sky130_fd_sc_hd__mux2_1 _12347_ (.A0(_05187_),
    .A1(\regs[11][10] ),
    .S(_06194_),
    .X(_06195_));
 sky130_fd_sc_hd__clkbuf_1 _12348_ (.A(_06195_),
    .X(_00649_));
 sky130_fd_sc_hd__mux2_1 _12349_ (.A0(_05224_),
    .A1(\regs[11][11] ),
    .S(_06194_),
    .X(_06196_));
 sky130_fd_sc_hd__clkbuf_1 _12350_ (.A(_06196_),
    .X(_00650_));
 sky130_fd_sc_hd__mux2_1 _12351_ (.A0(_05263_),
    .A1(\regs[11][12] ),
    .S(_06194_),
    .X(_06197_));
 sky130_fd_sc_hd__clkbuf_1 _12352_ (.A(_06197_),
    .X(_00651_));
 sky130_fd_sc_hd__mux2_1 _12353_ (.A0(_05296_),
    .A1(\regs[11][13] ),
    .S(_06194_),
    .X(_06198_));
 sky130_fd_sc_hd__clkbuf_1 _12354_ (.A(_06198_),
    .X(_00652_));
 sky130_fd_sc_hd__mux2_1 _12355_ (.A0(_05329_),
    .A1(\regs[11][14] ),
    .S(_06194_),
    .X(_06199_));
 sky130_fd_sc_hd__clkbuf_1 _12356_ (.A(_06199_),
    .X(_00653_));
 sky130_fd_sc_hd__mux2_1 _12357_ (.A0(_05359_),
    .A1(\regs[11][15] ),
    .S(_06194_),
    .X(_06200_));
 sky130_fd_sc_hd__clkbuf_1 _12358_ (.A(_06200_),
    .X(_00654_));
 sky130_fd_sc_hd__mux2_1 _12359_ (.A0(_05400_),
    .A1(\regs[11][16] ),
    .S(_06194_),
    .X(_06201_));
 sky130_fd_sc_hd__clkbuf_1 _12360_ (.A(_06201_),
    .X(_00655_));
 sky130_fd_sc_hd__mux2_1 _12361_ (.A0(_05424_),
    .A1(\regs[11][17] ),
    .S(_06194_),
    .X(_06202_));
 sky130_fd_sc_hd__clkbuf_1 _12362_ (.A(_06202_),
    .X(_00656_));
 sky130_fd_sc_hd__mux2_1 _12363_ (.A0(_05452_),
    .A1(\regs[11][18] ),
    .S(_06194_),
    .X(_06203_));
 sky130_fd_sc_hd__clkbuf_1 _12364_ (.A(_06203_),
    .X(_00657_));
 sky130_fd_sc_hd__mux2_1 _12365_ (.A0(_05477_),
    .A1(\regs[11][19] ),
    .S(_06194_),
    .X(_06204_));
 sky130_fd_sc_hd__clkbuf_1 _12366_ (.A(_06204_),
    .X(_00658_));
 sky130_fd_sc_hd__buf_8 _12367_ (.A(_06182_),
    .X(_06205_));
 sky130_fd_sc_hd__mux2_1 _12368_ (.A0(_05514_),
    .A1(\regs[11][20] ),
    .S(_06205_),
    .X(_06206_));
 sky130_fd_sc_hd__clkbuf_1 _12369_ (.A(_06206_),
    .X(_00659_));
 sky130_fd_sc_hd__mux2_1 _12370_ (.A0(_05541_),
    .A1(\regs[11][21] ),
    .S(_06205_),
    .X(_06207_));
 sky130_fd_sc_hd__clkbuf_1 _12371_ (.A(_06207_),
    .X(_00660_));
 sky130_fd_sc_hd__mux2_1 _12372_ (.A0(_05570_),
    .A1(\regs[11][22] ),
    .S(_06205_),
    .X(_06208_));
 sky130_fd_sc_hd__clkbuf_1 _12373_ (.A(_06208_),
    .X(_00661_));
 sky130_fd_sc_hd__mux2_1 _12374_ (.A0(_05600_),
    .A1(\regs[11][23] ),
    .S(_06205_),
    .X(_06209_));
 sky130_fd_sc_hd__clkbuf_1 _12375_ (.A(_06209_),
    .X(_00662_));
 sky130_fd_sc_hd__mux2_1 _12376_ (.A0(_05636_),
    .A1(\regs[11][24] ),
    .S(_06205_),
    .X(_06210_));
 sky130_fd_sc_hd__clkbuf_1 _12377_ (.A(_06210_),
    .X(_00663_));
 sky130_fd_sc_hd__mux2_1 _12378_ (.A0(_05660_),
    .A1(\regs[11][25] ),
    .S(_06205_),
    .X(_06211_));
 sky130_fd_sc_hd__clkbuf_1 _12379_ (.A(_06211_),
    .X(_00664_));
 sky130_fd_sc_hd__mux2_1 _12380_ (.A0(_05684_),
    .A1(\regs[11][26] ),
    .S(_06205_),
    .X(_06212_));
 sky130_fd_sc_hd__clkbuf_1 _12381_ (.A(_06212_),
    .X(_00665_));
 sky130_fd_sc_hd__mux2_1 _12382_ (.A0(_05708_),
    .A1(\regs[11][27] ),
    .S(_06205_),
    .X(_06213_));
 sky130_fd_sc_hd__clkbuf_1 _12383_ (.A(_06213_),
    .X(_00666_));
 sky130_fd_sc_hd__mux2_1 _12384_ (.A0(_05735_),
    .A1(\regs[11][28] ),
    .S(_06205_),
    .X(_06214_));
 sky130_fd_sc_hd__clkbuf_1 _12385_ (.A(_06214_),
    .X(_00667_));
 sky130_fd_sc_hd__mux2_1 _12386_ (.A0(_05763_),
    .A1(\regs[11][29] ),
    .S(_06205_),
    .X(_06215_));
 sky130_fd_sc_hd__clkbuf_1 _12387_ (.A(_06215_),
    .X(_00668_));
 sky130_fd_sc_hd__mux2_1 _12388_ (.A0(_05787_),
    .A1(\regs[11][30] ),
    .S(_06182_),
    .X(_06216_));
 sky130_fd_sc_hd__clkbuf_1 _12389_ (.A(_06216_),
    .X(_00669_));
 sky130_fd_sc_hd__mux2_1 _12390_ (.A0(_05811_),
    .A1(\regs[11][31] ),
    .S(_06182_),
    .X(_06217_));
 sky130_fd_sc_hd__clkbuf_1 _12391_ (.A(_06217_),
    .X(_00670_));
 sky130_fd_sc_hd__nand4_4 _12392_ (.A(_02313_),
    .B(_02315_),
    .C(_02241_),
    .D(_04765_),
    .Y(_06218_));
 sky130_fd_sc_hd__nor2_2 _12393_ (.A(_05958_),
    .B(_06218_),
    .Y(_06219_));
 sky130_fd_sc_hd__buf_6 _12394_ (.A(_06219_),
    .X(_06220_));
 sky130_fd_sc_hd__mux2_1 _12395_ (.A0(\regs[31][0] ),
    .A1(_05813_),
    .S(_06220_),
    .X(_06221_));
 sky130_fd_sc_hd__clkbuf_1 _12396_ (.A(_06221_),
    .X(_00671_));
 sky130_fd_sc_hd__mux2_1 _12397_ (.A0(\regs[31][1] ),
    .A1(_05819_),
    .S(_06220_),
    .X(_06222_));
 sky130_fd_sc_hd__clkbuf_1 _12398_ (.A(_06222_),
    .X(_00672_));
 sky130_fd_sc_hd__mux2_1 _12399_ (.A0(\regs[31][2] ),
    .A1(_05821_),
    .S(_06220_),
    .X(_06223_));
 sky130_fd_sc_hd__clkbuf_1 _12400_ (.A(_06223_),
    .X(_00673_));
 sky130_fd_sc_hd__mux2_1 _12401_ (.A0(\regs[31][3] ),
    .A1(_05823_),
    .S(_06220_),
    .X(_06224_));
 sky130_fd_sc_hd__clkbuf_1 _12402_ (.A(_06224_),
    .X(_00674_));
 sky130_fd_sc_hd__mux2_1 _12403_ (.A0(\regs[31][4] ),
    .A1(_05825_),
    .S(_06220_),
    .X(_06225_));
 sky130_fd_sc_hd__clkbuf_1 _12404_ (.A(_06225_),
    .X(_00675_));
 sky130_fd_sc_hd__mux2_1 _12405_ (.A0(\regs[31][5] ),
    .A1(_05827_),
    .S(_06220_),
    .X(_06226_));
 sky130_fd_sc_hd__clkbuf_1 _12406_ (.A(_06226_),
    .X(_00676_));
 sky130_fd_sc_hd__mux2_1 _12407_ (.A0(\regs[31][6] ),
    .A1(_05829_),
    .S(_06220_),
    .X(_06227_));
 sky130_fd_sc_hd__clkbuf_1 _12408_ (.A(_06227_),
    .X(_00677_));
 sky130_fd_sc_hd__mux2_1 _12409_ (.A0(\regs[31][7] ),
    .A1(_05831_),
    .S(_06220_),
    .X(_06228_));
 sky130_fd_sc_hd__clkbuf_1 _12410_ (.A(_06228_),
    .X(_00678_));
 sky130_fd_sc_hd__mux2_1 _12411_ (.A0(\regs[31][8] ),
    .A1(_05833_),
    .S(_06220_),
    .X(_06229_));
 sky130_fd_sc_hd__clkbuf_1 _12412_ (.A(_06229_),
    .X(_00679_));
 sky130_fd_sc_hd__mux2_1 _12413_ (.A0(\regs[31][9] ),
    .A1(_05835_),
    .S(_06220_),
    .X(_06230_));
 sky130_fd_sc_hd__clkbuf_1 _12414_ (.A(_06230_),
    .X(_00680_));
 sky130_fd_sc_hd__buf_4 _12415_ (.A(_06219_),
    .X(_06231_));
 sky130_fd_sc_hd__mux2_1 _12416_ (.A0(\regs[31][10] ),
    .A1(_05837_),
    .S(_06231_),
    .X(_06232_));
 sky130_fd_sc_hd__clkbuf_1 _12417_ (.A(_06232_),
    .X(_00681_));
 sky130_fd_sc_hd__mux2_1 _12418_ (.A0(\regs[31][11] ),
    .A1(_05840_),
    .S(_06231_),
    .X(_06233_));
 sky130_fd_sc_hd__clkbuf_1 _12419_ (.A(_06233_),
    .X(_00682_));
 sky130_fd_sc_hd__mux2_1 _12420_ (.A0(\regs[31][12] ),
    .A1(_05842_),
    .S(_06231_),
    .X(_06234_));
 sky130_fd_sc_hd__clkbuf_1 _12421_ (.A(_06234_),
    .X(_00683_));
 sky130_fd_sc_hd__mux2_1 _12422_ (.A0(\regs[31][13] ),
    .A1(_05844_),
    .S(_06231_),
    .X(_06235_));
 sky130_fd_sc_hd__clkbuf_1 _12423_ (.A(_06235_),
    .X(_00684_));
 sky130_fd_sc_hd__mux2_1 _12424_ (.A0(\regs[31][14] ),
    .A1(_05846_),
    .S(_06231_),
    .X(_06236_));
 sky130_fd_sc_hd__clkbuf_1 _12425_ (.A(_06236_),
    .X(_00685_));
 sky130_fd_sc_hd__mux2_1 _12426_ (.A0(\regs[31][15] ),
    .A1(_05848_),
    .S(_06231_),
    .X(_06237_));
 sky130_fd_sc_hd__clkbuf_1 _12427_ (.A(_06237_),
    .X(_00686_));
 sky130_fd_sc_hd__mux2_1 _12428_ (.A0(\regs[31][16] ),
    .A1(_05850_),
    .S(_06231_),
    .X(_06238_));
 sky130_fd_sc_hd__clkbuf_1 _12429_ (.A(_06238_),
    .X(_00687_));
 sky130_fd_sc_hd__mux2_1 _12430_ (.A0(\regs[31][17] ),
    .A1(_05852_),
    .S(_06231_),
    .X(_06239_));
 sky130_fd_sc_hd__clkbuf_1 _12431_ (.A(_06239_),
    .X(_00688_));
 sky130_fd_sc_hd__mux2_1 _12432_ (.A0(\regs[31][18] ),
    .A1(_05854_),
    .S(_06231_),
    .X(_06240_));
 sky130_fd_sc_hd__clkbuf_1 _12433_ (.A(_06240_),
    .X(_00689_));
 sky130_fd_sc_hd__mux2_1 _12434_ (.A0(\regs[31][19] ),
    .A1(_05856_),
    .S(_06231_),
    .X(_06241_));
 sky130_fd_sc_hd__clkbuf_1 _12435_ (.A(_06241_),
    .X(_00690_));
 sky130_fd_sc_hd__buf_4 _12436_ (.A(_06219_),
    .X(_06242_));
 sky130_fd_sc_hd__mux2_1 _12437_ (.A0(\regs[31][20] ),
    .A1(_05858_),
    .S(_06242_),
    .X(_06243_));
 sky130_fd_sc_hd__clkbuf_1 _12438_ (.A(_06243_),
    .X(_00691_));
 sky130_fd_sc_hd__mux2_1 _12439_ (.A0(\regs[31][21] ),
    .A1(_05861_),
    .S(_06242_),
    .X(_06244_));
 sky130_fd_sc_hd__clkbuf_1 _12440_ (.A(_06244_),
    .X(_00692_));
 sky130_fd_sc_hd__mux2_1 _12441_ (.A0(\regs[31][22] ),
    .A1(_05863_),
    .S(_06242_),
    .X(_06245_));
 sky130_fd_sc_hd__clkbuf_1 _12442_ (.A(_06245_),
    .X(_00693_));
 sky130_fd_sc_hd__mux2_1 _12443_ (.A0(\regs[31][23] ),
    .A1(_05865_),
    .S(_06242_),
    .X(_06246_));
 sky130_fd_sc_hd__clkbuf_1 _12444_ (.A(_06246_),
    .X(_00694_));
 sky130_fd_sc_hd__mux2_1 _12445_ (.A0(\regs[31][24] ),
    .A1(_05867_),
    .S(_06242_),
    .X(_06247_));
 sky130_fd_sc_hd__clkbuf_1 _12446_ (.A(_06247_),
    .X(_00695_));
 sky130_fd_sc_hd__mux2_1 _12447_ (.A0(\regs[31][25] ),
    .A1(_05869_),
    .S(_06242_),
    .X(_06248_));
 sky130_fd_sc_hd__clkbuf_1 _12448_ (.A(_06248_),
    .X(_00696_));
 sky130_fd_sc_hd__mux2_1 _12449_ (.A0(\regs[31][26] ),
    .A1(_05871_),
    .S(_06242_),
    .X(_06249_));
 sky130_fd_sc_hd__clkbuf_1 _12450_ (.A(_06249_),
    .X(_00697_));
 sky130_fd_sc_hd__mux2_1 _12451_ (.A0(\regs[31][27] ),
    .A1(_05873_),
    .S(_06242_),
    .X(_06250_));
 sky130_fd_sc_hd__clkbuf_1 _12452_ (.A(_06250_),
    .X(_00698_));
 sky130_fd_sc_hd__mux2_1 _12453_ (.A0(\regs[31][28] ),
    .A1(_05875_),
    .S(_06242_),
    .X(_06251_));
 sky130_fd_sc_hd__clkbuf_1 _12454_ (.A(_06251_),
    .X(_00699_));
 sky130_fd_sc_hd__mux2_1 _12455_ (.A0(\regs[31][29] ),
    .A1(_05877_),
    .S(_06242_),
    .X(_06252_));
 sky130_fd_sc_hd__clkbuf_1 _12456_ (.A(_06252_),
    .X(_00700_));
 sky130_fd_sc_hd__mux2_1 _12457_ (.A0(\regs[31][30] ),
    .A1(_05879_),
    .S(_06219_),
    .X(_06253_));
 sky130_fd_sc_hd__clkbuf_1 _12458_ (.A(_06253_),
    .X(_00701_));
 sky130_fd_sc_hd__mux2_1 _12459_ (.A0(\regs[31][31] ),
    .A1(_05881_),
    .S(_06219_),
    .X(_06254_));
 sky130_fd_sc_hd__clkbuf_1 _12460_ (.A(_06254_),
    .X(_00702_));
 sky130_fd_sc_hd__nor2_2 _12461_ (.A(_06072_),
    .B(_06218_),
    .Y(_06255_));
 sky130_fd_sc_hd__buf_6 _12462_ (.A(_06255_),
    .X(_06256_));
 sky130_fd_sc_hd__mux2_1 _12463_ (.A0(\regs[29][0] ),
    .A1(_05813_),
    .S(_06256_),
    .X(_06257_));
 sky130_fd_sc_hd__clkbuf_1 _12464_ (.A(_06257_),
    .X(_00703_));
 sky130_fd_sc_hd__mux2_1 _12465_ (.A0(\regs[29][1] ),
    .A1(_05819_),
    .S(_06256_),
    .X(_06258_));
 sky130_fd_sc_hd__clkbuf_1 _12466_ (.A(_06258_),
    .X(_00704_));
 sky130_fd_sc_hd__mux2_1 _12467_ (.A0(\regs[29][2] ),
    .A1(_05821_),
    .S(_06256_),
    .X(_06259_));
 sky130_fd_sc_hd__clkbuf_1 _12468_ (.A(_06259_),
    .X(_00705_));
 sky130_fd_sc_hd__mux2_1 _12469_ (.A0(\regs[29][3] ),
    .A1(_05823_),
    .S(_06256_),
    .X(_06260_));
 sky130_fd_sc_hd__clkbuf_1 _12470_ (.A(_06260_),
    .X(_00706_));
 sky130_fd_sc_hd__mux2_1 _12471_ (.A0(\regs[29][4] ),
    .A1(_05825_),
    .S(_06256_),
    .X(_06261_));
 sky130_fd_sc_hd__clkbuf_1 _12472_ (.A(_06261_),
    .X(_00707_));
 sky130_fd_sc_hd__mux2_1 _12473_ (.A0(\regs[29][5] ),
    .A1(_05827_),
    .S(_06256_),
    .X(_06262_));
 sky130_fd_sc_hd__clkbuf_1 _12474_ (.A(_06262_),
    .X(_00708_));
 sky130_fd_sc_hd__mux2_1 _12475_ (.A0(\regs[29][6] ),
    .A1(_05829_),
    .S(_06256_),
    .X(_06263_));
 sky130_fd_sc_hd__clkbuf_1 _12476_ (.A(_06263_),
    .X(_00709_));
 sky130_fd_sc_hd__mux2_1 _12477_ (.A0(\regs[29][7] ),
    .A1(_05831_),
    .S(_06256_),
    .X(_06264_));
 sky130_fd_sc_hd__clkbuf_1 _12478_ (.A(_06264_),
    .X(_00710_));
 sky130_fd_sc_hd__mux2_1 _12479_ (.A0(\regs[29][8] ),
    .A1(_05833_),
    .S(_06256_),
    .X(_06265_));
 sky130_fd_sc_hd__clkbuf_1 _12480_ (.A(_06265_),
    .X(_00711_));
 sky130_fd_sc_hd__mux2_1 _12481_ (.A0(\regs[29][9] ),
    .A1(_05835_),
    .S(_06256_),
    .X(_06266_));
 sky130_fd_sc_hd__clkbuf_1 _12482_ (.A(_06266_),
    .X(_00712_));
 sky130_fd_sc_hd__buf_6 _12483_ (.A(_06255_),
    .X(_06267_));
 sky130_fd_sc_hd__mux2_1 _12484_ (.A0(\regs[29][10] ),
    .A1(_05837_),
    .S(_06267_),
    .X(_06268_));
 sky130_fd_sc_hd__clkbuf_1 _12485_ (.A(_06268_),
    .X(_00713_));
 sky130_fd_sc_hd__mux2_1 _12486_ (.A0(\regs[29][11] ),
    .A1(_05840_),
    .S(_06267_),
    .X(_06269_));
 sky130_fd_sc_hd__clkbuf_1 _12487_ (.A(_06269_),
    .X(_00714_));
 sky130_fd_sc_hd__mux2_1 _12488_ (.A0(\regs[29][12] ),
    .A1(_05842_),
    .S(_06267_),
    .X(_06270_));
 sky130_fd_sc_hd__clkbuf_1 _12489_ (.A(_06270_),
    .X(_00715_));
 sky130_fd_sc_hd__mux2_1 _12490_ (.A0(\regs[29][13] ),
    .A1(_05844_),
    .S(_06267_),
    .X(_06271_));
 sky130_fd_sc_hd__clkbuf_1 _12491_ (.A(_06271_),
    .X(_00716_));
 sky130_fd_sc_hd__mux2_1 _12492_ (.A0(\regs[29][14] ),
    .A1(_05846_),
    .S(_06267_),
    .X(_06272_));
 sky130_fd_sc_hd__clkbuf_1 _12493_ (.A(_06272_),
    .X(_00717_));
 sky130_fd_sc_hd__mux2_1 _12494_ (.A0(\regs[29][15] ),
    .A1(_05848_),
    .S(_06267_),
    .X(_06273_));
 sky130_fd_sc_hd__clkbuf_1 _12495_ (.A(_06273_),
    .X(_00718_));
 sky130_fd_sc_hd__mux2_1 _12496_ (.A0(\regs[29][16] ),
    .A1(_05850_),
    .S(_06267_),
    .X(_06274_));
 sky130_fd_sc_hd__clkbuf_1 _12497_ (.A(_06274_),
    .X(_00719_));
 sky130_fd_sc_hd__mux2_1 _12498_ (.A0(\regs[29][17] ),
    .A1(_05852_),
    .S(_06267_),
    .X(_06275_));
 sky130_fd_sc_hd__clkbuf_1 _12499_ (.A(_06275_),
    .X(_00720_));
 sky130_fd_sc_hd__mux2_1 _12500_ (.A0(\regs[29][18] ),
    .A1(_05854_),
    .S(_06267_),
    .X(_06276_));
 sky130_fd_sc_hd__clkbuf_1 _12501_ (.A(_06276_),
    .X(_00721_));
 sky130_fd_sc_hd__mux2_1 _12502_ (.A0(\regs[29][19] ),
    .A1(_05856_),
    .S(_06267_),
    .X(_06277_));
 sky130_fd_sc_hd__clkbuf_1 _12503_ (.A(_06277_),
    .X(_00722_));
 sky130_fd_sc_hd__buf_4 _12504_ (.A(_06255_),
    .X(_06278_));
 sky130_fd_sc_hd__mux2_1 _12505_ (.A0(\regs[29][20] ),
    .A1(_05858_),
    .S(_06278_),
    .X(_06279_));
 sky130_fd_sc_hd__clkbuf_1 _12506_ (.A(_06279_),
    .X(_00723_));
 sky130_fd_sc_hd__mux2_1 _12507_ (.A0(\regs[29][21] ),
    .A1(_05861_),
    .S(_06278_),
    .X(_06280_));
 sky130_fd_sc_hd__clkbuf_1 _12508_ (.A(_06280_),
    .X(_00724_));
 sky130_fd_sc_hd__mux2_1 _12509_ (.A0(\regs[29][22] ),
    .A1(_05863_),
    .S(_06278_),
    .X(_06281_));
 sky130_fd_sc_hd__clkbuf_1 _12510_ (.A(_06281_),
    .X(_00725_));
 sky130_fd_sc_hd__mux2_1 _12511_ (.A0(\regs[29][23] ),
    .A1(_05865_),
    .S(_06278_),
    .X(_06282_));
 sky130_fd_sc_hd__clkbuf_1 _12512_ (.A(_06282_),
    .X(_00726_));
 sky130_fd_sc_hd__mux2_1 _12513_ (.A0(\regs[29][24] ),
    .A1(_05867_),
    .S(_06278_),
    .X(_06283_));
 sky130_fd_sc_hd__clkbuf_1 _12514_ (.A(_06283_),
    .X(_00727_));
 sky130_fd_sc_hd__mux2_1 _12515_ (.A0(\regs[29][25] ),
    .A1(_05869_),
    .S(_06278_),
    .X(_06284_));
 sky130_fd_sc_hd__clkbuf_1 _12516_ (.A(_06284_),
    .X(_00728_));
 sky130_fd_sc_hd__mux2_1 _12517_ (.A0(\regs[29][26] ),
    .A1(_05871_),
    .S(_06278_),
    .X(_06285_));
 sky130_fd_sc_hd__clkbuf_1 _12518_ (.A(_06285_),
    .X(_00729_));
 sky130_fd_sc_hd__mux2_1 _12519_ (.A0(\regs[29][27] ),
    .A1(_05873_),
    .S(_06278_),
    .X(_06286_));
 sky130_fd_sc_hd__clkbuf_1 _12520_ (.A(_06286_),
    .X(_00730_));
 sky130_fd_sc_hd__mux2_1 _12521_ (.A0(\regs[29][28] ),
    .A1(_05875_),
    .S(_06278_),
    .X(_06287_));
 sky130_fd_sc_hd__clkbuf_1 _12522_ (.A(_06287_),
    .X(_00731_));
 sky130_fd_sc_hd__mux2_1 _12523_ (.A0(\regs[29][29] ),
    .A1(_05877_),
    .S(_06278_),
    .X(_06288_));
 sky130_fd_sc_hd__clkbuf_1 _12524_ (.A(_06288_),
    .X(_00732_));
 sky130_fd_sc_hd__mux2_1 _12525_ (.A0(\regs[29][30] ),
    .A1(_05879_),
    .S(_06255_),
    .X(_06289_));
 sky130_fd_sc_hd__clkbuf_1 _12526_ (.A(_06289_),
    .X(_00733_));
 sky130_fd_sc_hd__mux2_1 _12527_ (.A0(\regs[29][31] ),
    .A1(_05881_),
    .S(_06255_),
    .X(_06290_));
 sky130_fd_sc_hd__clkbuf_1 _12528_ (.A(_06290_),
    .X(_00734_));
 sky130_fd_sc_hd__buf_2 _12529_ (.A(_04761_),
    .X(_06291_));
 sky130_fd_sc_hd__nor2_4 _12530_ (.A(_04757_),
    .B(_05958_),
    .Y(_06292_));
 sky130_fd_sc_hd__buf_6 _12531_ (.A(_06292_),
    .X(_06293_));
 sky130_fd_sc_hd__mux2_1 _12532_ (.A0(\regs[3][0] ),
    .A1(_06291_),
    .S(_06293_),
    .X(_06294_));
 sky130_fd_sc_hd__clkbuf_1 _12533_ (.A(_06294_),
    .X(_00735_));
 sky130_fd_sc_hd__buf_2 _12534_ (.A(_04817_),
    .X(_06295_));
 sky130_fd_sc_hd__mux2_1 _12535_ (.A0(\regs[3][1] ),
    .A1(_06295_),
    .S(_06293_),
    .X(_06296_));
 sky130_fd_sc_hd__clkbuf_1 _12536_ (.A(_06296_),
    .X(_00736_));
 sky130_fd_sc_hd__buf_2 _12537_ (.A(_04857_),
    .X(_06297_));
 sky130_fd_sc_hd__mux2_1 _12538_ (.A0(\regs[3][2] ),
    .A1(_06297_),
    .S(_06293_),
    .X(_06298_));
 sky130_fd_sc_hd__clkbuf_1 _12539_ (.A(_06298_),
    .X(_00737_));
 sky130_fd_sc_hd__buf_2 _12540_ (.A(_04903_),
    .X(_06299_));
 sky130_fd_sc_hd__mux2_1 _12541_ (.A0(\regs[3][3] ),
    .A1(_06299_),
    .S(_06293_),
    .X(_06300_));
 sky130_fd_sc_hd__clkbuf_1 _12542_ (.A(_06300_),
    .X(_00738_));
 sky130_fd_sc_hd__buf_2 _12543_ (.A(_04951_),
    .X(_06301_));
 sky130_fd_sc_hd__mux2_1 _12544_ (.A0(\regs[3][4] ),
    .A1(_06301_),
    .S(_06293_),
    .X(_06302_));
 sky130_fd_sc_hd__clkbuf_1 _12545_ (.A(_06302_),
    .X(_00739_));
 sky130_fd_sc_hd__buf_2 _12546_ (.A(_04991_),
    .X(_06303_));
 sky130_fd_sc_hd__mux2_1 _12547_ (.A0(\regs[3][5] ),
    .A1(_06303_),
    .S(_06293_),
    .X(_06304_));
 sky130_fd_sc_hd__clkbuf_1 _12548_ (.A(_06304_),
    .X(_00740_));
 sky130_fd_sc_hd__buf_2 _12549_ (.A(_05029_),
    .X(_06305_));
 sky130_fd_sc_hd__mux2_1 _12550_ (.A0(\regs[3][6] ),
    .A1(_06305_),
    .S(_06293_),
    .X(_06306_));
 sky130_fd_sc_hd__clkbuf_1 _12551_ (.A(_06306_),
    .X(_00741_));
 sky130_fd_sc_hd__buf_2 _12552_ (.A(_05079_),
    .X(_06307_));
 sky130_fd_sc_hd__mux2_1 _12553_ (.A0(\regs[3][7] ),
    .A1(_06307_),
    .S(_06293_),
    .X(_06308_));
 sky130_fd_sc_hd__clkbuf_1 _12554_ (.A(_06308_),
    .X(_00742_));
 sky130_fd_sc_hd__buf_2 _12555_ (.A(_05120_),
    .X(_06309_));
 sky130_fd_sc_hd__mux2_1 _12556_ (.A0(\regs[3][8] ),
    .A1(_06309_),
    .S(_06293_),
    .X(_06310_));
 sky130_fd_sc_hd__clkbuf_1 _12557_ (.A(_06310_),
    .X(_00743_));
 sky130_fd_sc_hd__buf_2 _12558_ (.A(_05156_),
    .X(_06311_));
 sky130_fd_sc_hd__mux2_1 _12559_ (.A0(\regs[3][9] ),
    .A1(_06311_),
    .S(_06293_),
    .X(_06312_));
 sky130_fd_sc_hd__clkbuf_1 _12560_ (.A(_06312_),
    .X(_00744_));
 sky130_fd_sc_hd__clkbuf_4 _12561_ (.A(_05186_),
    .X(_06313_));
 sky130_fd_sc_hd__clkbuf_8 _12562_ (.A(_06292_),
    .X(_06314_));
 sky130_fd_sc_hd__mux2_1 _12563_ (.A0(\regs[3][10] ),
    .A1(_06313_),
    .S(_06314_),
    .X(_06315_));
 sky130_fd_sc_hd__clkbuf_1 _12564_ (.A(_06315_),
    .X(_00745_));
 sky130_fd_sc_hd__clkbuf_4 _12565_ (.A(_05223_),
    .X(_06316_));
 sky130_fd_sc_hd__mux2_1 _12566_ (.A0(\regs[3][11] ),
    .A1(_06316_),
    .S(_06314_),
    .X(_06317_));
 sky130_fd_sc_hd__clkbuf_1 _12567_ (.A(_06317_),
    .X(_00746_));
 sky130_fd_sc_hd__clkbuf_4 _12568_ (.A(_05262_),
    .X(_06318_));
 sky130_fd_sc_hd__mux2_1 _12569_ (.A0(\regs[3][12] ),
    .A1(_06318_),
    .S(_06314_),
    .X(_06319_));
 sky130_fd_sc_hd__clkbuf_1 _12570_ (.A(_06319_),
    .X(_00747_));
 sky130_fd_sc_hd__buf_2 _12571_ (.A(_05295_),
    .X(_06320_));
 sky130_fd_sc_hd__mux2_1 _12572_ (.A0(\regs[3][13] ),
    .A1(_06320_),
    .S(_06314_),
    .X(_06321_));
 sky130_fd_sc_hd__clkbuf_1 _12573_ (.A(_06321_),
    .X(_00748_));
 sky130_fd_sc_hd__clkbuf_4 _12574_ (.A(_05328_),
    .X(_06322_));
 sky130_fd_sc_hd__mux2_1 _12575_ (.A0(\regs[3][14] ),
    .A1(_06322_),
    .S(_06314_),
    .X(_06323_));
 sky130_fd_sc_hd__clkbuf_1 _12576_ (.A(_06323_),
    .X(_00749_));
 sky130_fd_sc_hd__buf_2 _12577_ (.A(_05358_),
    .X(_06324_));
 sky130_fd_sc_hd__mux2_1 _12578_ (.A0(\regs[3][15] ),
    .A1(_06324_),
    .S(_06314_),
    .X(_06325_));
 sky130_fd_sc_hd__clkbuf_1 _12579_ (.A(_06325_),
    .X(_00750_));
 sky130_fd_sc_hd__clkbuf_4 _12580_ (.A(_05399_),
    .X(_06326_));
 sky130_fd_sc_hd__mux2_1 _12581_ (.A0(\regs[3][16] ),
    .A1(_06326_),
    .S(_06314_),
    .X(_06327_));
 sky130_fd_sc_hd__clkbuf_1 _12582_ (.A(_06327_),
    .X(_00751_));
 sky130_fd_sc_hd__clkbuf_4 _12583_ (.A(_05423_),
    .X(_06328_));
 sky130_fd_sc_hd__mux2_1 _12584_ (.A0(\regs[3][17] ),
    .A1(_06328_),
    .S(_06314_),
    .X(_06329_));
 sky130_fd_sc_hd__clkbuf_1 _12585_ (.A(_06329_),
    .X(_00752_));
 sky130_fd_sc_hd__clkbuf_4 _12586_ (.A(_05451_),
    .X(_06330_));
 sky130_fd_sc_hd__mux2_1 _12587_ (.A0(\regs[3][18] ),
    .A1(_06330_),
    .S(_06314_),
    .X(_06331_));
 sky130_fd_sc_hd__clkbuf_1 _12588_ (.A(_06331_),
    .X(_00753_));
 sky130_fd_sc_hd__clkbuf_4 _12589_ (.A(_05476_),
    .X(_06332_));
 sky130_fd_sc_hd__mux2_1 _12590_ (.A0(\regs[3][19] ),
    .A1(_06332_),
    .S(_06314_),
    .X(_06333_));
 sky130_fd_sc_hd__clkbuf_1 _12591_ (.A(_06333_),
    .X(_00754_));
 sky130_fd_sc_hd__buf_2 _12592_ (.A(_05513_),
    .X(_06334_));
 sky130_fd_sc_hd__buf_6 _12593_ (.A(_06292_),
    .X(_06335_));
 sky130_fd_sc_hd__mux2_1 _12594_ (.A0(\regs[3][20] ),
    .A1(_06334_),
    .S(_06335_),
    .X(_06336_));
 sky130_fd_sc_hd__clkbuf_1 _12595_ (.A(_06336_),
    .X(_00755_));
 sky130_fd_sc_hd__buf_4 _12596_ (.A(_05540_),
    .X(_06337_));
 sky130_fd_sc_hd__mux2_1 _12597_ (.A0(\regs[3][21] ),
    .A1(_06337_),
    .S(_06335_),
    .X(_06338_));
 sky130_fd_sc_hd__clkbuf_1 _12598_ (.A(_06338_),
    .X(_00756_));
 sky130_fd_sc_hd__clkbuf_4 _12599_ (.A(_05569_),
    .X(_06339_));
 sky130_fd_sc_hd__mux2_1 _12600_ (.A0(\regs[3][22] ),
    .A1(_06339_),
    .S(_06335_),
    .X(_06340_));
 sky130_fd_sc_hd__clkbuf_1 _12601_ (.A(_06340_),
    .X(_00757_));
 sky130_fd_sc_hd__buf_2 _12602_ (.A(_05599_),
    .X(_06341_));
 sky130_fd_sc_hd__mux2_1 _12603_ (.A0(\regs[3][23] ),
    .A1(_06341_),
    .S(_06335_),
    .X(_06342_));
 sky130_fd_sc_hd__clkbuf_1 _12604_ (.A(_06342_),
    .X(_00758_));
 sky130_fd_sc_hd__buf_2 _12605_ (.A(_05635_),
    .X(_06343_));
 sky130_fd_sc_hd__mux2_1 _12606_ (.A0(\regs[3][24] ),
    .A1(_06343_),
    .S(_06335_),
    .X(_06344_));
 sky130_fd_sc_hd__clkbuf_1 _12607_ (.A(_06344_),
    .X(_00759_));
 sky130_fd_sc_hd__buf_2 _12608_ (.A(_05659_),
    .X(_06345_));
 sky130_fd_sc_hd__mux2_1 _12609_ (.A0(\regs[3][25] ),
    .A1(_06345_),
    .S(_06335_),
    .X(_06346_));
 sky130_fd_sc_hd__clkbuf_1 _12610_ (.A(_06346_),
    .X(_00760_));
 sky130_fd_sc_hd__clkbuf_4 _12611_ (.A(_05683_),
    .X(_06347_));
 sky130_fd_sc_hd__mux2_1 _12612_ (.A0(\regs[3][26] ),
    .A1(_06347_),
    .S(_06335_),
    .X(_06348_));
 sky130_fd_sc_hd__clkbuf_1 _12613_ (.A(_06348_),
    .X(_00761_));
 sky130_fd_sc_hd__clkbuf_4 _12614_ (.A(_05707_),
    .X(_06349_));
 sky130_fd_sc_hd__mux2_1 _12615_ (.A0(\regs[3][27] ),
    .A1(_06349_),
    .S(_06335_),
    .X(_06350_));
 sky130_fd_sc_hd__clkbuf_1 _12616_ (.A(_06350_),
    .X(_00762_));
 sky130_fd_sc_hd__buf_2 _12617_ (.A(_05734_),
    .X(_06351_));
 sky130_fd_sc_hd__mux2_1 _12618_ (.A0(\regs[3][28] ),
    .A1(_06351_),
    .S(_06335_),
    .X(_06352_));
 sky130_fd_sc_hd__clkbuf_1 _12619_ (.A(_06352_),
    .X(_00763_));
 sky130_fd_sc_hd__clkbuf_4 _12620_ (.A(_05762_),
    .X(_06353_));
 sky130_fd_sc_hd__mux2_1 _12621_ (.A0(\regs[3][29] ),
    .A1(_06353_),
    .S(_06335_),
    .X(_06354_));
 sky130_fd_sc_hd__clkbuf_1 _12622_ (.A(_06354_),
    .X(_00764_));
 sky130_fd_sc_hd__buf_2 _12623_ (.A(_05786_),
    .X(_06355_));
 sky130_fd_sc_hd__mux2_1 _12624_ (.A0(\regs[3][30] ),
    .A1(_06355_),
    .S(_06292_),
    .X(_06356_));
 sky130_fd_sc_hd__clkbuf_1 _12625_ (.A(_06356_),
    .X(_00765_));
 sky130_fd_sc_hd__buf_2 _12626_ (.A(_05810_),
    .X(_06357_));
 sky130_fd_sc_hd__mux2_1 _12627_ (.A0(\regs[3][31] ),
    .A1(_06357_),
    .S(_06292_),
    .X(_06358_));
 sky130_fd_sc_hd__clkbuf_1 _12628_ (.A(_06358_),
    .X(_00766_));
 sky130_fd_sc_hd__nor2_4 _12629_ (.A(_05958_),
    .B(_06145_),
    .Y(_06359_));
 sky130_fd_sc_hd__buf_6 _12630_ (.A(_06359_),
    .X(_06360_));
 sky130_fd_sc_hd__mux2_1 _12631_ (.A0(\regs[19][0] ),
    .A1(_06291_),
    .S(_06360_),
    .X(_06361_));
 sky130_fd_sc_hd__clkbuf_1 _12632_ (.A(_06361_),
    .X(_00767_));
 sky130_fd_sc_hd__mux2_1 _12633_ (.A0(\regs[19][1] ),
    .A1(_06295_),
    .S(_06360_),
    .X(_06362_));
 sky130_fd_sc_hd__clkbuf_1 _12634_ (.A(_06362_),
    .X(_00768_));
 sky130_fd_sc_hd__mux2_1 _12635_ (.A0(\regs[19][2] ),
    .A1(_06297_),
    .S(_06360_),
    .X(_06363_));
 sky130_fd_sc_hd__clkbuf_1 _12636_ (.A(_06363_),
    .X(_00769_));
 sky130_fd_sc_hd__mux2_1 _12637_ (.A0(\regs[19][3] ),
    .A1(_06299_),
    .S(_06360_),
    .X(_06364_));
 sky130_fd_sc_hd__clkbuf_1 _12638_ (.A(_06364_),
    .X(_00770_));
 sky130_fd_sc_hd__mux2_1 _12639_ (.A0(\regs[19][4] ),
    .A1(_06301_),
    .S(_06360_),
    .X(_06365_));
 sky130_fd_sc_hd__clkbuf_1 _12640_ (.A(_06365_),
    .X(_00771_));
 sky130_fd_sc_hd__mux2_1 _12641_ (.A0(\regs[19][5] ),
    .A1(_06303_),
    .S(_06360_),
    .X(_06366_));
 sky130_fd_sc_hd__clkbuf_1 _12642_ (.A(_06366_),
    .X(_00772_));
 sky130_fd_sc_hd__mux2_1 _12643_ (.A0(\regs[19][6] ),
    .A1(_06305_),
    .S(_06360_),
    .X(_06367_));
 sky130_fd_sc_hd__clkbuf_1 _12644_ (.A(_06367_),
    .X(_00773_));
 sky130_fd_sc_hd__mux2_1 _12645_ (.A0(\regs[19][7] ),
    .A1(_06307_),
    .S(_06360_),
    .X(_06368_));
 sky130_fd_sc_hd__clkbuf_1 _12646_ (.A(_06368_),
    .X(_00774_));
 sky130_fd_sc_hd__mux2_1 _12647_ (.A0(\regs[19][8] ),
    .A1(_06309_),
    .S(_06360_),
    .X(_06369_));
 sky130_fd_sc_hd__clkbuf_1 _12648_ (.A(_06369_),
    .X(_00775_));
 sky130_fd_sc_hd__mux2_1 _12649_ (.A0(\regs[19][9] ),
    .A1(_06311_),
    .S(_06360_),
    .X(_06370_));
 sky130_fd_sc_hd__clkbuf_1 _12650_ (.A(_06370_),
    .X(_00776_));
 sky130_fd_sc_hd__clkbuf_8 _12651_ (.A(_06359_),
    .X(_06371_));
 sky130_fd_sc_hd__mux2_1 _12652_ (.A0(\regs[19][10] ),
    .A1(_06313_),
    .S(_06371_),
    .X(_06372_));
 sky130_fd_sc_hd__clkbuf_1 _12653_ (.A(_06372_),
    .X(_00777_));
 sky130_fd_sc_hd__mux2_1 _12654_ (.A0(\regs[19][11] ),
    .A1(_06316_),
    .S(_06371_),
    .X(_06373_));
 sky130_fd_sc_hd__clkbuf_1 _12655_ (.A(_06373_),
    .X(_00778_));
 sky130_fd_sc_hd__mux2_1 _12656_ (.A0(\regs[19][12] ),
    .A1(_06318_),
    .S(_06371_),
    .X(_06374_));
 sky130_fd_sc_hd__clkbuf_1 _12657_ (.A(_06374_),
    .X(_00779_));
 sky130_fd_sc_hd__mux2_1 _12658_ (.A0(\regs[19][13] ),
    .A1(_06320_),
    .S(_06371_),
    .X(_06375_));
 sky130_fd_sc_hd__clkbuf_1 _12659_ (.A(_06375_),
    .X(_00780_));
 sky130_fd_sc_hd__mux2_1 _12660_ (.A0(\regs[19][14] ),
    .A1(_06322_),
    .S(_06371_),
    .X(_06376_));
 sky130_fd_sc_hd__clkbuf_1 _12661_ (.A(_06376_),
    .X(_00781_));
 sky130_fd_sc_hd__mux2_1 _12662_ (.A0(\regs[19][15] ),
    .A1(_06324_),
    .S(_06371_),
    .X(_06377_));
 sky130_fd_sc_hd__clkbuf_1 _12663_ (.A(_06377_),
    .X(_00782_));
 sky130_fd_sc_hd__mux2_1 _12664_ (.A0(\regs[19][16] ),
    .A1(_06326_),
    .S(_06371_),
    .X(_06378_));
 sky130_fd_sc_hd__clkbuf_1 _12665_ (.A(_06378_),
    .X(_00783_));
 sky130_fd_sc_hd__mux2_1 _12666_ (.A0(\regs[19][17] ),
    .A1(_06328_),
    .S(_06371_),
    .X(_06379_));
 sky130_fd_sc_hd__clkbuf_1 _12667_ (.A(_06379_),
    .X(_00784_));
 sky130_fd_sc_hd__mux2_1 _12668_ (.A0(\regs[19][18] ),
    .A1(_06330_),
    .S(_06371_),
    .X(_06380_));
 sky130_fd_sc_hd__clkbuf_1 _12669_ (.A(_06380_),
    .X(_00785_));
 sky130_fd_sc_hd__mux2_1 _12670_ (.A0(\regs[19][19] ),
    .A1(_06332_),
    .S(_06371_),
    .X(_06381_));
 sky130_fd_sc_hd__clkbuf_1 _12671_ (.A(_06381_),
    .X(_00786_));
 sky130_fd_sc_hd__buf_6 _12672_ (.A(_06359_),
    .X(_06382_));
 sky130_fd_sc_hd__mux2_1 _12673_ (.A0(\regs[19][20] ),
    .A1(_06334_),
    .S(_06382_),
    .X(_06383_));
 sky130_fd_sc_hd__clkbuf_1 _12674_ (.A(_06383_),
    .X(_00787_));
 sky130_fd_sc_hd__mux2_1 _12675_ (.A0(\regs[19][21] ),
    .A1(_06337_),
    .S(_06382_),
    .X(_06384_));
 sky130_fd_sc_hd__clkbuf_1 _12676_ (.A(_06384_),
    .X(_00788_));
 sky130_fd_sc_hd__mux2_1 _12677_ (.A0(\regs[19][22] ),
    .A1(_06339_),
    .S(_06382_),
    .X(_06385_));
 sky130_fd_sc_hd__clkbuf_1 _12678_ (.A(_06385_),
    .X(_00789_));
 sky130_fd_sc_hd__mux2_1 _12679_ (.A0(\regs[19][23] ),
    .A1(_06341_),
    .S(_06382_),
    .X(_06386_));
 sky130_fd_sc_hd__clkbuf_1 _12680_ (.A(_06386_),
    .X(_00790_));
 sky130_fd_sc_hd__mux2_1 _12681_ (.A0(\regs[19][24] ),
    .A1(_06343_),
    .S(_06382_),
    .X(_06387_));
 sky130_fd_sc_hd__clkbuf_1 _12682_ (.A(_06387_),
    .X(_00791_));
 sky130_fd_sc_hd__mux2_1 _12683_ (.A0(\regs[19][25] ),
    .A1(_06345_),
    .S(_06382_),
    .X(_06388_));
 sky130_fd_sc_hd__clkbuf_1 _12684_ (.A(_06388_),
    .X(_00792_));
 sky130_fd_sc_hd__mux2_1 _12685_ (.A0(\regs[19][26] ),
    .A1(_06347_),
    .S(_06382_),
    .X(_06389_));
 sky130_fd_sc_hd__clkbuf_1 _12686_ (.A(_06389_),
    .X(_00793_));
 sky130_fd_sc_hd__mux2_1 _12687_ (.A0(\regs[19][27] ),
    .A1(_06349_),
    .S(_06382_),
    .X(_06390_));
 sky130_fd_sc_hd__clkbuf_1 _12688_ (.A(_06390_),
    .X(_00794_));
 sky130_fd_sc_hd__mux2_1 _12689_ (.A0(\regs[19][28] ),
    .A1(_06351_),
    .S(_06382_),
    .X(_06391_));
 sky130_fd_sc_hd__clkbuf_1 _12690_ (.A(_06391_),
    .X(_00795_));
 sky130_fd_sc_hd__mux2_1 _12691_ (.A0(\regs[19][29] ),
    .A1(_06353_),
    .S(_06382_),
    .X(_06392_));
 sky130_fd_sc_hd__clkbuf_1 _12692_ (.A(_06392_),
    .X(_00796_));
 sky130_fd_sc_hd__mux2_1 _12693_ (.A0(\regs[19][30] ),
    .A1(_06355_),
    .S(_06359_),
    .X(_06393_));
 sky130_fd_sc_hd__clkbuf_1 _12694_ (.A(_06393_),
    .X(_00797_));
 sky130_fd_sc_hd__mux2_1 _12695_ (.A0(\regs[19][31] ),
    .A1(_06357_),
    .S(_06359_),
    .X(_06394_));
 sky130_fd_sc_hd__clkbuf_1 _12696_ (.A(_06394_),
    .X(_00798_));
 sky130_fd_sc_hd__nand2_4 _12697_ (.A(_06031_),
    .B(_05815_),
    .Y(_06395_));
 sky130_fd_sc_hd__buf_6 _12698_ (.A(_06395_),
    .X(_06396_));
 sky130_fd_sc_hd__mux2_1 _12699_ (.A0(_04762_),
    .A1(\regs[4][0] ),
    .S(_06396_),
    .X(_06397_));
 sky130_fd_sc_hd__clkbuf_1 _12700_ (.A(_06397_),
    .X(_00799_));
 sky130_fd_sc_hd__mux2_1 _12701_ (.A0(_04818_),
    .A1(\regs[4][1] ),
    .S(_06396_),
    .X(_06398_));
 sky130_fd_sc_hd__clkbuf_1 _12702_ (.A(_06398_),
    .X(_00800_));
 sky130_fd_sc_hd__mux2_1 _12703_ (.A0(_04858_),
    .A1(\regs[4][2] ),
    .S(_06396_),
    .X(_06399_));
 sky130_fd_sc_hd__clkbuf_1 _12704_ (.A(_06399_),
    .X(_00801_));
 sky130_fd_sc_hd__mux2_1 _12705_ (.A0(_04904_),
    .A1(\regs[4][3] ),
    .S(_06396_),
    .X(_06400_));
 sky130_fd_sc_hd__clkbuf_1 _12706_ (.A(_06400_),
    .X(_00802_));
 sky130_fd_sc_hd__mux2_1 _12707_ (.A0(_04952_),
    .A1(\regs[4][4] ),
    .S(_06396_),
    .X(_06401_));
 sky130_fd_sc_hd__clkbuf_1 _12708_ (.A(_06401_),
    .X(_00803_));
 sky130_fd_sc_hd__mux2_1 _12709_ (.A0(_04992_),
    .A1(\regs[4][5] ),
    .S(_06396_),
    .X(_06402_));
 sky130_fd_sc_hd__clkbuf_1 _12710_ (.A(_06402_),
    .X(_00804_));
 sky130_fd_sc_hd__mux2_1 _12711_ (.A0(_05030_),
    .A1(\regs[4][6] ),
    .S(_06396_),
    .X(_06403_));
 sky130_fd_sc_hd__clkbuf_1 _12712_ (.A(_06403_),
    .X(_00805_));
 sky130_fd_sc_hd__mux2_1 _12713_ (.A0(_05080_),
    .A1(\regs[4][7] ),
    .S(_06396_),
    .X(_06404_));
 sky130_fd_sc_hd__clkbuf_1 _12714_ (.A(_06404_),
    .X(_00806_));
 sky130_fd_sc_hd__mux2_1 _12715_ (.A0(_05121_),
    .A1(\regs[4][8] ),
    .S(_06396_),
    .X(_06405_));
 sky130_fd_sc_hd__clkbuf_1 _12716_ (.A(_06405_),
    .X(_00807_));
 sky130_fd_sc_hd__mux2_1 _12717_ (.A0(_05157_),
    .A1(\regs[4][9] ),
    .S(_06396_),
    .X(_06406_));
 sky130_fd_sc_hd__clkbuf_1 _12718_ (.A(_06406_),
    .X(_00808_));
 sky130_fd_sc_hd__buf_4 _12719_ (.A(_06395_),
    .X(_06407_));
 sky130_fd_sc_hd__mux2_1 _12720_ (.A0(_05187_),
    .A1(\regs[4][10] ),
    .S(_06407_),
    .X(_06408_));
 sky130_fd_sc_hd__clkbuf_1 _12721_ (.A(_06408_),
    .X(_00809_));
 sky130_fd_sc_hd__mux2_1 _12722_ (.A0(_05224_),
    .A1(\regs[4][11] ),
    .S(_06407_),
    .X(_06409_));
 sky130_fd_sc_hd__clkbuf_1 _12723_ (.A(_06409_),
    .X(_00810_));
 sky130_fd_sc_hd__mux2_1 _12724_ (.A0(_05263_),
    .A1(\regs[4][12] ),
    .S(_06407_),
    .X(_06410_));
 sky130_fd_sc_hd__clkbuf_1 _12725_ (.A(_06410_),
    .X(_00811_));
 sky130_fd_sc_hd__mux2_1 _12726_ (.A0(_05296_),
    .A1(\regs[4][13] ),
    .S(_06407_),
    .X(_06411_));
 sky130_fd_sc_hd__clkbuf_1 _12727_ (.A(_06411_),
    .X(_00812_));
 sky130_fd_sc_hd__mux2_1 _12728_ (.A0(_05329_),
    .A1(\regs[4][14] ),
    .S(_06407_),
    .X(_06412_));
 sky130_fd_sc_hd__clkbuf_1 _12729_ (.A(_06412_),
    .X(_00813_));
 sky130_fd_sc_hd__mux2_1 _12730_ (.A0(_05359_),
    .A1(\regs[4][15] ),
    .S(_06407_),
    .X(_06413_));
 sky130_fd_sc_hd__clkbuf_1 _12731_ (.A(_06413_),
    .X(_00814_));
 sky130_fd_sc_hd__mux2_1 _12732_ (.A0(_05400_),
    .A1(\regs[4][16] ),
    .S(_06407_),
    .X(_06414_));
 sky130_fd_sc_hd__clkbuf_1 _12733_ (.A(_06414_),
    .X(_00815_));
 sky130_fd_sc_hd__mux2_1 _12734_ (.A0(_05424_),
    .A1(\regs[4][17] ),
    .S(_06407_),
    .X(_06415_));
 sky130_fd_sc_hd__clkbuf_1 _12735_ (.A(_06415_),
    .X(_00816_));
 sky130_fd_sc_hd__mux2_1 _12736_ (.A0(_05452_),
    .A1(\regs[4][18] ),
    .S(_06407_),
    .X(_06416_));
 sky130_fd_sc_hd__clkbuf_1 _12737_ (.A(_06416_),
    .X(_00817_));
 sky130_fd_sc_hd__mux2_1 _12738_ (.A0(_05477_),
    .A1(\regs[4][19] ),
    .S(_06407_),
    .X(_06417_));
 sky130_fd_sc_hd__clkbuf_1 _12739_ (.A(_06417_),
    .X(_00818_));
 sky130_fd_sc_hd__buf_8 _12740_ (.A(_06395_),
    .X(_06418_));
 sky130_fd_sc_hd__mux2_1 _12741_ (.A0(_05514_),
    .A1(\regs[4][20] ),
    .S(_06418_),
    .X(_06419_));
 sky130_fd_sc_hd__clkbuf_1 _12742_ (.A(_06419_),
    .X(_00819_));
 sky130_fd_sc_hd__mux2_1 _12743_ (.A0(_05541_),
    .A1(\regs[4][21] ),
    .S(_06418_),
    .X(_06420_));
 sky130_fd_sc_hd__clkbuf_1 _12744_ (.A(_06420_),
    .X(_00820_));
 sky130_fd_sc_hd__mux2_1 _12745_ (.A0(_05570_),
    .A1(\regs[4][22] ),
    .S(_06418_),
    .X(_06421_));
 sky130_fd_sc_hd__clkbuf_1 _12746_ (.A(_06421_),
    .X(_00821_));
 sky130_fd_sc_hd__mux2_1 _12747_ (.A0(_05600_),
    .A1(\regs[4][23] ),
    .S(_06418_),
    .X(_06422_));
 sky130_fd_sc_hd__clkbuf_1 _12748_ (.A(_06422_),
    .X(_00822_));
 sky130_fd_sc_hd__mux2_1 _12749_ (.A0(_05636_),
    .A1(\regs[4][24] ),
    .S(_06418_),
    .X(_06423_));
 sky130_fd_sc_hd__clkbuf_1 _12750_ (.A(_06423_),
    .X(_00823_));
 sky130_fd_sc_hd__mux2_1 _12751_ (.A0(_05660_),
    .A1(\regs[4][25] ),
    .S(_06418_),
    .X(_06424_));
 sky130_fd_sc_hd__clkbuf_1 _12752_ (.A(_06424_),
    .X(_00824_));
 sky130_fd_sc_hd__mux2_1 _12753_ (.A0(_05684_),
    .A1(\regs[4][26] ),
    .S(_06418_),
    .X(_06425_));
 sky130_fd_sc_hd__clkbuf_1 _12754_ (.A(_06425_),
    .X(_00825_));
 sky130_fd_sc_hd__mux2_1 _12755_ (.A0(_05708_),
    .A1(\regs[4][27] ),
    .S(_06418_),
    .X(_06426_));
 sky130_fd_sc_hd__clkbuf_1 _12756_ (.A(_06426_),
    .X(_00826_));
 sky130_fd_sc_hd__mux2_1 _12757_ (.A0(_05735_),
    .A1(\regs[4][28] ),
    .S(_06418_),
    .X(_06427_));
 sky130_fd_sc_hd__clkbuf_1 _12758_ (.A(_06427_),
    .X(_00827_));
 sky130_fd_sc_hd__mux2_1 _12759_ (.A0(_05763_),
    .A1(\regs[4][29] ),
    .S(_06418_),
    .X(_06428_));
 sky130_fd_sc_hd__clkbuf_1 _12760_ (.A(_06428_),
    .X(_00828_));
 sky130_fd_sc_hd__mux2_1 _12761_ (.A0(_05787_),
    .A1(\regs[4][30] ),
    .S(_06395_),
    .X(_06429_));
 sky130_fd_sc_hd__clkbuf_1 _12762_ (.A(_06429_),
    .X(_00829_));
 sky130_fd_sc_hd__mux2_1 _12763_ (.A0(_05811_),
    .A1(\regs[4][31] ),
    .S(_06395_),
    .X(_06430_));
 sky130_fd_sc_hd__clkbuf_1 _12764_ (.A(_06430_),
    .X(_00830_));
 sky130_fd_sc_hd__inv_2 _12765_ (.A(_06070_),
    .Y(_00072_));
 sky130_fd_sc_hd__and2_1 _12766_ (.A(_00068_),
    .B(\regs[0][0] ),
    .X(_06431_));
 sky130_fd_sc_hd__clkbuf_1 _12767_ (.A(_06431_),
    .X(_00832_));
 sky130_fd_sc_hd__and2_1 _12768_ (.A(_00068_),
    .B(\regs[0][1] ),
    .X(_06432_));
 sky130_fd_sc_hd__clkbuf_1 _12769_ (.A(_06432_),
    .X(_00833_));
 sky130_fd_sc_hd__and2_1 _12770_ (.A(_00068_),
    .B(\regs[0][2] ),
    .X(_06433_));
 sky130_fd_sc_hd__clkbuf_1 _12771_ (.A(_06433_),
    .X(_00834_));
 sky130_fd_sc_hd__and2_1 _12772_ (.A(_00068_),
    .B(\regs[0][3] ),
    .X(_06434_));
 sky130_fd_sc_hd__clkbuf_1 _12773_ (.A(_06434_),
    .X(_00835_));
 sky130_fd_sc_hd__and2_1 _12774_ (.A(_00068_),
    .B(\regs[0][4] ),
    .X(_06435_));
 sky130_fd_sc_hd__clkbuf_1 _12775_ (.A(_06435_),
    .X(_00836_));
 sky130_fd_sc_hd__and2_1 _12776_ (.A(_00068_),
    .B(\regs[0][5] ),
    .X(_06436_));
 sky130_fd_sc_hd__clkbuf_1 _12777_ (.A(_06436_),
    .X(_00837_));
 sky130_fd_sc_hd__and2_1 _12778_ (.A(_00068_),
    .B(\regs[0][6] ),
    .X(_06437_));
 sky130_fd_sc_hd__clkbuf_1 _12779_ (.A(_06437_),
    .X(_00838_));
 sky130_fd_sc_hd__and2_1 _12780_ (.A(_00068_),
    .B(\regs[0][7] ),
    .X(_06438_));
 sky130_fd_sc_hd__clkbuf_1 _12781_ (.A(_06438_),
    .X(_00839_));
 sky130_fd_sc_hd__and2_1 _12782_ (.A(_00068_),
    .B(\regs[0][8] ),
    .X(_06439_));
 sky130_fd_sc_hd__clkbuf_1 _12783_ (.A(_06439_),
    .X(_00840_));
 sky130_fd_sc_hd__buf_4 _12784_ (.A(_06068_),
    .X(_06440_));
 sky130_fd_sc_hd__and2_1 _12785_ (.A(_06440_),
    .B(\regs[0][9] ),
    .X(_06441_));
 sky130_fd_sc_hd__clkbuf_1 _12786_ (.A(_06441_),
    .X(_00841_));
 sky130_fd_sc_hd__and2_1 _12787_ (.A(_06440_),
    .B(\regs[0][10] ),
    .X(_06442_));
 sky130_fd_sc_hd__clkbuf_1 _12788_ (.A(_06442_),
    .X(_00842_));
 sky130_fd_sc_hd__and2_1 _12789_ (.A(_06440_),
    .B(\regs[0][11] ),
    .X(_06443_));
 sky130_fd_sc_hd__clkbuf_1 _12790_ (.A(_06443_),
    .X(_00843_));
 sky130_fd_sc_hd__and2_1 _12791_ (.A(_06440_),
    .B(\regs[0][12] ),
    .X(_06444_));
 sky130_fd_sc_hd__clkbuf_1 _12792_ (.A(_06444_),
    .X(_00844_));
 sky130_fd_sc_hd__and2_1 _12793_ (.A(_06440_),
    .B(\regs[0][13] ),
    .X(_06445_));
 sky130_fd_sc_hd__clkbuf_1 _12794_ (.A(_06445_),
    .X(_00845_));
 sky130_fd_sc_hd__and2_1 _12795_ (.A(_06440_),
    .B(\regs[0][14] ),
    .X(_06446_));
 sky130_fd_sc_hd__clkbuf_1 _12796_ (.A(_06446_),
    .X(_00846_));
 sky130_fd_sc_hd__and2_1 _12797_ (.A(_06440_),
    .B(\regs[0][15] ),
    .X(_06447_));
 sky130_fd_sc_hd__clkbuf_1 _12798_ (.A(_06447_),
    .X(_00847_));
 sky130_fd_sc_hd__and2_1 _12799_ (.A(_06440_),
    .B(\regs[0][16] ),
    .X(_06448_));
 sky130_fd_sc_hd__clkbuf_1 _12800_ (.A(_06448_),
    .X(_00848_));
 sky130_fd_sc_hd__and2_1 _12801_ (.A(_06440_),
    .B(\regs[0][17] ),
    .X(_06449_));
 sky130_fd_sc_hd__clkbuf_1 _12802_ (.A(_06449_),
    .X(_00849_));
 sky130_fd_sc_hd__and2_1 _12803_ (.A(_06440_),
    .B(\regs[0][18] ),
    .X(_06450_));
 sky130_fd_sc_hd__clkbuf_1 _12804_ (.A(_06450_),
    .X(_00850_));
 sky130_fd_sc_hd__buf_4 _12805_ (.A(_06068_),
    .X(_06451_));
 sky130_fd_sc_hd__and2_1 _12806_ (.A(_06451_),
    .B(\regs[0][19] ),
    .X(_06452_));
 sky130_fd_sc_hd__clkbuf_1 _12807_ (.A(_06452_),
    .X(_00851_));
 sky130_fd_sc_hd__and2_1 _12808_ (.A(_06451_),
    .B(\regs[0][20] ),
    .X(_06453_));
 sky130_fd_sc_hd__clkbuf_1 _12809_ (.A(_06453_),
    .X(_00852_));
 sky130_fd_sc_hd__and2_1 _12810_ (.A(_06451_),
    .B(\regs[0][21] ),
    .X(_06454_));
 sky130_fd_sc_hd__clkbuf_1 _12811_ (.A(_06454_),
    .X(_00853_));
 sky130_fd_sc_hd__and2_1 _12812_ (.A(_06451_),
    .B(\regs[0][22] ),
    .X(_06455_));
 sky130_fd_sc_hd__clkbuf_1 _12813_ (.A(_06455_),
    .X(_00854_));
 sky130_fd_sc_hd__and2_1 _12814_ (.A(_06451_),
    .B(\regs[0][23] ),
    .X(_06456_));
 sky130_fd_sc_hd__clkbuf_1 _12815_ (.A(_06456_),
    .X(_00855_));
 sky130_fd_sc_hd__and2_1 _12816_ (.A(_06451_),
    .B(\regs[0][24] ),
    .X(_06457_));
 sky130_fd_sc_hd__clkbuf_1 _12817_ (.A(_06457_),
    .X(_00856_));
 sky130_fd_sc_hd__and2_1 _12818_ (.A(_06451_),
    .B(\regs[0][25] ),
    .X(_06458_));
 sky130_fd_sc_hd__clkbuf_1 _12819_ (.A(_06458_),
    .X(_00857_));
 sky130_fd_sc_hd__and2_1 _12820_ (.A(_06451_),
    .B(\regs[0][26] ),
    .X(_06459_));
 sky130_fd_sc_hd__clkbuf_1 _12821_ (.A(_06459_),
    .X(_00858_));
 sky130_fd_sc_hd__and2_1 _12822_ (.A(_06451_),
    .B(\regs[0][27] ),
    .X(_06460_));
 sky130_fd_sc_hd__clkbuf_1 _12823_ (.A(_06460_),
    .X(_00859_));
 sky130_fd_sc_hd__and2_1 _12824_ (.A(_06451_),
    .B(\regs[0][28] ),
    .X(_06461_));
 sky130_fd_sc_hd__clkbuf_1 _12825_ (.A(_06461_),
    .X(_00860_));
 sky130_fd_sc_hd__and2_1 _12826_ (.A(_06068_),
    .B(\regs[0][29] ),
    .X(_06462_));
 sky130_fd_sc_hd__clkbuf_1 _12827_ (.A(_06462_),
    .X(_00861_));
 sky130_fd_sc_hd__and2_1 _12828_ (.A(_06068_),
    .B(\regs[0][30] ),
    .X(_06463_));
 sky130_fd_sc_hd__clkbuf_1 _12829_ (.A(_06463_),
    .X(_00862_));
 sky130_fd_sc_hd__and2_1 _12830_ (.A(_06068_),
    .B(\regs[0][31] ),
    .X(_06464_));
 sky130_fd_sc_hd__clkbuf_1 _12831_ (.A(_06464_),
    .X(_00863_));
 sky130_fd_sc_hd__nor2_4 _12832_ (.A(_05883_),
    .B(_06145_),
    .Y(_06465_));
 sky130_fd_sc_hd__buf_6 _12833_ (.A(_06465_),
    .X(_06466_));
 sky130_fd_sc_hd__mux2_1 _12834_ (.A0(\regs[18][0] ),
    .A1(_06291_),
    .S(_06466_),
    .X(_06467_));
 sky130_fd_sc_hd__clkbuf_1 _12835_ (.A(_06467_),
    .X(_00864_));
 sky130_fd_sc_hd__mux2_1 _12836_ (.A0(\regs[18][1] ),
    .A1(_06295_),
    .S(_06466_),
    .X(_06468_));
 sky130_fd_sc_hd__clkbuf_1 _12837_ (.A(_06468_),
    .X(_00865_));
 sky130_fd_sc_hd__mux2_1 _12838_ (.A0(\regs[18][2] ),
    .A1(_06297_),
    .S(_06466_),
    .X(_06469_));
 sky130_fd_sc_hd__clkbuf_1 _12839_ (.A(_06469_),
    .X(_00866_));
 sky130_fd_sc_hd__mux2_1 _12840_ (.A0(\regs[18][3] ),
    .A1(_06299_),
    .S(_06466_),
    .X(_06470_));
 sky130_fd_sc_hd__clkbuf_1 _12841_ (.A(_06470_),
    .X(_00867_));
 sky130_fd_sc_hd__mux2_1 _12842_ (.A0(\regs[18][4] ),
    .A1(_06301_),
    .S(_06466_),
    .X(_06471_));
 sky130_fd_sc_hd__clkbuf_1 _12843_ (.A(_06471_),
    .X(_00868_));
 sky130_fd_sc_hd__mux2_1 _12844_ (.A0(\regs[18][5] ),
    .A1(_06303_),
    .S(_06466_),
    .X(_06472_));
 sky130_fd_sc_hd__clkbuf_1 _12845_ (.A(_06472_),
    .X(_00869_));
 sky130_fd_sc_hd__mux2_1 _12846_ (.A0(\regs[18][6] ),
    .A1(_06305_),
    .S(_06466_),
    .X(_06473_));
 sky130_fd_sc_hd__clkbuf_1 _12847_ (.A(_06473_),
    .X(_00870_));
 sky130_fd_sc_hd__mux2_1 _12848_ (.A0(\regs[18][7] ),
    .A1(_06307_),
    .S(_06466_),
    .X(_06474_));
 sky130_fd_sc_hd__clkbuf_1 _12849_ (.A(_06474_),
    .X(_00871_));
 sky130_fd_sc_hd__mux2_1 _12850_ (.A0(\regs[18][8] ),
    .A1(_06309_),
    .S(_06466_),
    .X(_06475_));
 sky130_fd_sc_hd__clkbuf_1 _12851_ (.A(_06475_),
    .X(_00872_));
 sky130_fd_sc_hd__mux2_1 _12852_ (.A0(\regs[18][9] ),
    .A1(_06311_),
    .S(_06466_),
    .X(_06476_));
 sky130_fd_sc_hd__clkbuf_1 _12853_ (.A(_06476_),
    .X(_00873_));
 sky130_fd_sc_hd__buf_6 _12854_ (.A(_06465_),
    .X(_06477_));
 sky130_fd_sc_hd__mux2_1 _12855_ (.A0(\regs[18][10] ),
    .A1(_06313_),
    .S(_06477_),
    .X(_06478_));
 sky130_fd_sc_hd__clkbuf_1 _12856_ (.A(_06478_),
    .X(_00874_));
 sky130_fd_sc_hd__mux2_1 _12857_ (.A0(\regs[18][11] ),
    .A1(_06316_),
    .S(_06477_),
    .X(_06479_));
 sky130_fd_sc_hd__clkbuf_1 _12858_ (.A(_06479_),
    .X(_00875_));
 sky130_fd_sc_hd__mux2_1 _12859_ (.A0(\regs[18][12] ),
    .A1(_06318_),
    .S(_06477_),
    .X(_06480_));
 sky130_fd_sc_hd__clkbuf_1 _12860_ (.A(_06480_),
    .X(_00876_));
 sky130_fd_sc_hd__mux2_1 _12861_ (.A0(\regs[18][13] ),
    .A1(_06320_),
    .S(_06477_),
    .X(_06481_));
 sky130_fd_sc_hd__clkbuf_1 _12862_ (.A(_06481_),
    .X(_00877_));
 sky130_fd_sc_hd__mux2_1 _12863_ (.A0(\regs[18][14] ),
    .A1(_06322_),
    .S(_06477_),
    .X(_06482_));
 sky130_fd_sc_hd__clkbuf_1 _12864_ (.A(_06482_),
    .X(_00878_));
 sky130_fd_sc_hd__mux2_1 _12865_ (.A0(\regs[18][15] ),
    .A1(_06324_),
    .S(_06477_),
    .X(_06483_));
 sky130_fd_sc_hd__clkbuf_1 _12866_ (.A(_06483_),
    .X(_00879_));
 sky130_fd_sc_hd__mux2_1 _12867_ (.A0(\regs[18][16] ),
    .A1(_06326_),
    .S(_06477_),
    .X(_06484_));
 sky130_fd_sc_hd__clkbuf_1 _12868_ (.A(_06484_),
    .X(_00880_));
 sky130_fd_sc_hd__mux2_1 _12869_ (.A0(\regs[18][17] ),
    .A1(_06328_),
    .S(_06477_),
    .X(_06485_));
 sky130_fd_sc_hd__clkbuf_1 _12870_ (.A(_06485_),
    .X(_00881_));
 sky130_fd_sc_hd__mux2_1 _12871_ (.A0(\regs[18][18] ),
    .A1(_06330_),
    .S(_06477_),
    .X(_06486_));
 sky130_fd_sc_hd__clkbuf_1 _12872_ (.A(_06486_),
    .X(_00882_));
 sky130_fd_sc_hd__mux2_1 _12873_ (.A0(\regs[18][19] ),
    .A1(_06332_),
    .S(_06477_),
    .X(_06487_));
 sky130_fd_sc_hd__clkbuf_1 _12874_ (.A(_06487_),
    .X(_00883_));
 sky130_fd_sc_hd__buf_6 _12875_ (.A(_06465_),
    .X(_06488_));
 sky130_fd_sc_hd__mux2_1 _12876_ (.A0(\regs[18][20] ),
    .A1(_06334_),
    .S(_06488_),
    .X(_06489_));
 sky130_fd_sc_hd__clkbuf_1 _12877_ (.A(_06489_),
    .X(_00884_));
 sky130_fd_sc_hd__mux2_1 _12878_ (.A0(\regs[18][21] ),
    .A1(_06337_),
    .S(_06488_),
    .X(_06490_));
 sky130_fd_sc_hd__clkbuf_1 _12879_ (.A(_06490_),
    .X(_00885_));
 sky130_fd_sc_hd__mux2_1 _12880_ (.A0(\regs[18][22] ),
    .A1(_06339_),
    .S(_06488_),
    .X(_06491_));
 sky130_fd_sc_hd__clkbuf_1 _12881_ (.A(_06491_),
    .X(_00886_));
 sky130_fd_sc_hd__mux2_1 _12882_ (.A0(\regs[18][23] ),
    .A1(_06341_),
    .S(_06488_),
    .X(_06492_));
 sky130_fd_sc_hd__clkbuf_1 _12883_ (.A(_06492_),
    .X(_00887_));
 sky130_fd_sc_hd__mux2_1 _12884_ (.A0(\regs[18][24] ),
    .A1(_06343_),
    .S(_06488_),
    .X(_06493_));
 sky130_fd_sc_hd__clkbuf_1 _12885_ (.A(_06493_),
    .X(_00888_));
 sky130_fd_sc_hd__mux2_1 _12886_ (.A0(\regs[18][25] ),
    .A1(_06345_),
    .S(_06488_),
    .X(_06494_));
 sky130_fd_sc_hd__clkbuf_1 _12887_ (.A(_06494_),
    .X(_00889_));
 sky130_fd_sc_hd__mux2_1 _12888_ (.A0(\regs[18][26] ),
    .A1(_06347_),
    .S(_06488_),
    .X(_06495_));
 sky130_fd_sc_hd__clkbuf_1 _12889_ (.A(_06495_),
    .X(_00890_));
 sky130_fd_sc_hd__mux2_1 _12890_ (.A0(\regs[18][27] ),
    .A1(_06349_),
    .S(_06488_),
    .X(_06496_));
 sky130_fd_sc_hd__clkbuf_1 _12891_ (.A(_06496_),
    .X(_00891_));
 sky130_fd_sc_hd__mux2_1 _12892_ (.A0(\regs[18][28] ),
    .A1(_06351_),
    .S(_06488_),
    .X(_06497_));
 sky130_fd_sc_hd__clkbuf_1 _12893_ (.A(_06497_),
    .X(_00892_));
 sky130_fd_sc_hd__mux2_1 _12894_ (.A0(\regs[18][29] ),
    .A1(_06353_),
    .S(_06488_),
    .X(_06498_));
 sky130_fd_sc_hd__clkbuf_1 _12895_ (.A(_06498_),
    .X(_00893_));
 sky130_fd_sc_hd__mux2_1 _12896_ (.A0(\regs[18][30] ),
    .A1(_06355_),
    .S(_06465_),
    .X(_06499_));
 sky130_fd_sc_hd__clkbuf_1 _12897_ (.A(_06499_),
    .X(_00894_));
 sky130_fd_sc_hd__mux2_1 _12898_ (.A0(\regs[18][31] ),
    .A1(_06357_),
    .S(_06465_),
    .X(_06500_));
 sky130_fd_sc_hd__clkbuf_1 _12899_ (.A(_06500_),
    .X(_00895_));
 sky130_fd_sc_hd__nor2_4 _12900_ (.A(_06072_),
    .B(_04757_),
    .Y(_06501_));
 sky130_fd_sc_hd__buf_6 _12901_ (.A(_06501_),
    .X(_06502_));
 sky130_fd_sc_hd__mux2_1 _12902_ (.A0(\regs[1][0] ),
    .A1(_06291_),
    .S(_06502_),
    .X(_06503_));
 sky130_fd_sc_hd__clkbuf_1 _12903_ (.A(_06503_),
    .X(_00896_));
 sky130_fd_sc_hd__mux2_1 _12904_ (.A0(\regs[1][1] ),
    .A1(_06295_),
    .S(_06502_),
    .X(_06504_));
 sky130_fd_sc_hd__clkbuf_1 _12905_ (.A(_06504_),
    .X(_00897_));
 sky130_fd_sc_hd__mux2_1 _12906_ (.A0(\regs[1][2] ),
    .A1(_06297_),
    .S(_06502_),
    .X(_06505_));
 sky130_fd_sc_hd__clkbuf_1 _12907_ (.A(_06505_),
    .X(_00898_));
 sky130_fd_sc_hd__mux2_1 _12908_ (.A0(\regs[1][3] ),
    .A1(_06299_),
    .S(_06502_),
    .X(_06506_));
 sky130_fd_sc_hd__clkbuf_1 _12909_ (.A(_06506_),
    .X(_00899_));
 sky130_fd_sc_hd__mux2_1 _12910_ (.A0(\regs[1][4] ),
    .A1(_06301_),
    .S(_06502_),
    .X(_06507_));
 sky130_fd_sc_hd__clkbuf_1 _12911_ (.A(_06507_),
    .X(_00900_));
 sky130_fd_sc_hd__mux2_1 _12912_ (.A0(\regs[1][5] ),
    .A1(_06303_),
    .S(_06502_),
    .X(_06508_));
 sky130_fd_sc_hd__clkbuf_1 _12913_ (.A(_06508_),
    .X(_00901_));
 sky130_fd_sc_hd__mux2_1 _12914_ (.A0(\regs[1][6] ),
    .A1(_06305_),
    .S(_06502_),
    .X(_06509_));
 sky130_fd_sc_hd__clkbuf_1 _12915_ (.A(_06509_),
    .X(_00902_));
 sky130_fd_sc_hd__mux2_1 _12916_ (.A0(\regs[1][7] ),
    .A1(_06307_),
    .S(_06502_),
    .X(_06510_));
 sky130_fd_sc_hd__clkbuf_1 _12917_ (.A(_06510_),
    .X(_00903_));
 sky130_fd_sc_hd__mux2_1 _12918_ (.A0(\regs[1][8] ),
    .A1(_06309_),
    .S(_06502_),
    .X(_06511_));
 sky130_fd_sc_hd__clkbuf_1 _12919_ (.A(_06511_),
    .X(_00904_));
 sky130_fd_sc_hd__mux2_1 _12920_ (.A0(\regs[1][9] ),
    .A1(_06311_),
    .S(_06502_),
    .X(_06512_));
 sky130_fd_sc_hd__clkbuf_1 _12921_ (.A(_06512_),
    .X(_00905_));
 sky130_fd_sc_hd__clkbuf_8 _12922_ (.A(_06501_),
    .X(_06513_));
 sky130_fd_sc_hd__mux2_1 _12923_ (.A0(\regs[1][10] ),
    .A1(_06313_),
    .S(_06513_),
    .X(_06514_));
 sky130_fd_sc_hd__clkbuf_1 _12924_ (.A(_06514_),
    .X(_00906_));
 sky130_fd_sc_hd__mux2_1 _12925_ (.A0(\regs[1][11] ),
    .A1(_06316_),
    .S(_06513_),
    .X(_06515_));
 sky130_fd_sc_hd__clkbuf_1 _12926_ (.A(_06515_),
    .X(_00907_));
 sky130_fd_sc_hd__mux2_1 _12927_ (.A0(\regs[1][12] ),
    .A1(_06318_),
    .S(_06513_),
    .X(_06516_));
 sky130_fd_sc_hd__clkbuf_1 _12928_ (.A(_06516_),
    .X(_00908_));
 sky130_fd_sc_hd__mux2_1 _12929_ (.A0(\regs[1][13] ),
    .A1(_06320_),
    .S(_06513_),
    .X(_06517_));
 sky130_fd_sc_hd__clkbuf_1 _12930_ (.A(_06517_),
    .X(_00909_));
 sky130_fd_sc_hd__mux2_1 _12931_ (.A0(\regs[1][14] ),
    .A1(_06322_),
    .S(_06513_),
    .X(_06518_));
 sky130_fd_sc_hd__clkbuf_1 _12932_ (.A(_06518_),
    .X(_00910_));
 sky130_fd_sc_hd__mux2_1 _12933_ (.A0(\regs[1][15] ),
    .A1(_06324_),
    .S(_06513_),
    .X(_06519_));
 sky130_fd_sc_hd__clkbuf_1 _12934_ (.A(_06519_),
    .X(_00911_));
 sky130_fd_sc_hd__mux2_1 _12935_ (.A0(\regs[1][16] ),
    .A1(_06326_),
    .S(_06513_),
    .X(_06520_));
 sky130_fd_sc_hd__clkbuf_1 _12936_ (.A(_06520_),
    .X(_00912_));
 sky130_fd_sc_hd__mux2_1 _12937_ (.A0(\regs[1][17] ),
    .A1(_06328_),
    .S(_06513_),
    .X(_06521_));
 sky130_fd_sc_hd__clkbuf_1 _12938_ (.A(_06521_),
    .X(_00913_));
 sky130_fd_sc_hd__mux2_1 _12939_ (.A0(\regs[1][18] ),
    .A1(_06330_),
    .S(_06513_),
    .X(_06522_));
 sky130_fd_sc_hd__clkbuf_1 _12940_ (.A(_06522_),
    .X(_00914_));
 sky130_fd_sc_hd__mux2_1 _12941_ (.A0(\regs[1][19] ),
    .A1(_06332_),
    .S(_06513_),
    .X(_06523_));
 sky130_fd_sc_hd__clkbuf_1 _12942_ (.A(_06523_),
    .X(_00915_));
 sky130_fd_sc_hd__buf_6 _12943_ (.A(_06501_),
    .X(_06524_));
 sky130_fd_sc_hd__mux2_1 _12944_ (.A0(\regs[1][20] ),
    .A1(_06334_),
    .S(_06524_),
    .X(_06525_));
 sky130_fd_sc_hd__clkbuf_1 _12945_ (.A(_06525_),
    .X(_00916_));
 sky130_fd_sc_hd__mux2_1 _12946_ (.A0(\regs[1][21] ),
    .A1(_06337_),
    .S(_06524_),
    .X(_06526_));
 sky130_fd_sc_hd__clkbuf_1 _12947_ (.A(_06526_),
    .X(_00917_));
 sky130_fd_sc_hd__mux2_1 _12948_ (.A0(\regs[1][22] ),
    .A1(_06339_),
    .S(_06524_),
    .X(_06527_));
 sky130_fd_sc_hd__clkbuf_1 _12949_ (.A(_06527_),
    .X(_00918_));
 sky130_fd_sc_hd__mux2_1 _12950_ (.A0(\regs[1][23] ),
    .A1(_06341_),
    .S(_06524_),
    .X(_06528_));
 sky130_fd_sc_hd__clkbuf_1 _12951_ (.A(_06528_),
    .X(_00919_));
 sky130_fd_sc_hd__mux2_1 _12952_ (.A0(\regs[1][24] ),
    .A1(_06343_),
    .S(_06524_),
    .X(_06529_));
 sky130_fd_sc_hd__clkbuf_1 _12953_ (.A(_06529_),
    .X(_00920_));
 sky130_fd_sc_hd__mux2_1 _12954_ (.A0(\regs[1][25] ),
    .A1(_06345_),
    .S(_06524_),
    .X(_06530_));
 sky130_fd_sc_hd__clkbuf_1 _12955_ (.A(_06530_),
    .X(_00921_));
 sky130_fd_sc_hd__mux2_1 _12956_ (.A0(\regs[1][26] ),
    .A1(_06347_),
    .S(_06524_),
    .X(_06531_));
 sky130_fd_sc_hd__clkbuf_1 _12957_ (.A(_06531_),
    .X(_00922_));
 sky130_fd_sc_hd__mux2_1 _12958_ (.A0(\regs[1][27] ),
    .A1(_06349_),
    .S(_06524_),
    .X(_06532_));
 sky130_fd_sc_hd__clkbuf_1 _12959_ (.A(_06532_),
    .X(_00923_));
 sky130_fd_sc_hd__mux2_1 _12960_ (.A0(\regs[1][28] ),
    .A1(_06351_),
    .S(_06524_),
    .X(_06533_));
 sky130_fd_sc_hd__clkbuf_1 _12961_ (.A(_06533_),
    .X(_00924_));
 sky130_fd_sc_hd__mux2_1 _12962_ (.A0(\regs[1][29] ),
    .A1(_06353_),
    .S(_06524_),
    .X(_06534_));
 sky130_fd_sc_hd__clkbuf_1 _12963_ (.A(_06534_),
    .X(_00925_));
 sky130_fd_sc_hd__mux2_1 _12964_ (.A0(\regs[1][30] ),
    .A1(_06355_),
    .S(_06501_),
    .X(_06535_));
 sky130_fd_sc_hd__clkbuf_1 _12965_ (.A(_06535_),
    .X(_00926_));
 sky130_fd_sc_hd__mux2_1 _12966_ (.A0(\regs[1][31] ),
    .A1(_06357_),
    .S(_06501_),
    .X(_06536_));
 sky130_fd_sc_hd__clkbuf_1 _12967_ (.A(_06536_),
    .X(_00927_));
 sky130_fd_sc_hd__nand4b_4 _12968_ (.A_N(_02315_),
    .B(_02241_),
    .C(_04765_),
    .D(_02313_),
    .Y(_06537_));
 sky130_fd_sc_hd__or2_4 _12969_ (.A(_04758_),
    .B(_06537_),
    .X(_06538_));
 sky130_fd_sc_hd__buf_6 _12970_ (.A(_06538_),
    .X(_06539_));
 sky130_fd_sc_hd__mux2_1 _12971_ (.A0(_04762_),
    .A1(\regs[20][0] ),
    .S(_06539_),
    .X(_06540_));
 sky130_fd_sc_hd__clkbuf_1 _12972_ (.A(_06540_),
    .X(_00928_));
 sky130_fd_sc_hd__mux2_1 _12973_ (.A0(_04818_),
    .A1(\regs[20][1] ),
    .S(_06539_),
    .X(_06541_));
 sky130_fd_sc_hd__clkbuf_1 _12974_ (.A(_06541_),
    .X(_00929_));
 sky130_fd_sc_hd__mux2_1 _12975_ (.A0(_04858_),
    .A1(\regs[20][2] ),
    .S(_06539_),
    .X(_06542_));
 sky130_fd_sc_hd__clkbuf_1 _12976_ (.A(_06542_),
    .X(_00930_));
 sky130_fd_sc_hd__mux2_1 _12977_ (.A0(_04904_),
    .A1(\regs[20][3] ),
    .S(_06539_),
    .X(_06543_));
 sky130_fd_sc_hd__clkbuf_1 _12978_ (.A(_06543_),
    .X(_00931_));
 sky130_fd_sc_hd__mux2_1 _12979_ (.A0(_04952_),
    .A1(\regs[20][4] ),
    .S(_06539_),
    .X(_06544_));
 sky130_fd_sc_hd__clkbuf_1 _12980_ (.A(_06544_),
    .X(_00932_));
 sky130_fd_sc_hd__mux2_1 _12981_ (.A0(_04992_),
    .A1(\regs[20][5] ),
    .S(_06539_),
    .X(_06545_));
 sky130_fd_sc_hd__clkbuf_1 _12982_ (.A(_06545_),
    .X(_00933_));
 sky130_fd_sc_hd__mux2_1 _12983_ (.A0(_05030_),
    .A1(\regs[20][6] ),
    .S(_06539_),
    .X(_06546_));
 sky130_fd_sc_hd__clkbuf_1 _12984_ (.A(_06546_),
    .X(_00934_));
 sky130_fd_sc_hd__mux2_1 _12985_ (.A0(_05080_),
    .A1(\regs[20][7] ),
    .S(_06539_),
    .X(_06547_));
 sky130_fd_sc_hd__clkbuf_1 _12986_ (.A(_06547_),
    .X(_00935_));
 sky130_fd_sc_hd__mux2_1 _12987_ (.A0(_05121_),
    .A1(\regs[20][8] ),
    .S(_06539_),
    .X(_06548_));
 sky130_fd_sc_hd__clkbuf_1 _12988_ (.A(_06548_),
    .X(_00936_));
 sky130_fd_sc_hd__mux2_1 _12989_ (.A0(_05157_),
    .A1(\regs[20][9] ),
    .S(_06539_),
    .X(_06549_));
 sky130_fd_sc_hd__clkbuf_1 _12990_ (.A(_06549_),
    .X(_00937_));
 sky130_fd_sc_hd__buf_6 _12991_ (.A(_06538_),
    .X(_06550_));
 sky130_fd_sc_hd__mux2_1 _12992_ (.A0(_05187_),
    .A1(\regs[20][10] ),
    .S(_06550_),
    .X(_06551_));
 sky130_fd_sc_hd__clkbuf_1 _12993_ (.A(_06551_),
    .X(_00938_));
 sky130_fd_sc_hd__mux2_1 _12994_ (.A0(_05224_),
    .A1(\regs[20][11] ),
    .S(_06550_),
    .X(_06552_));
 sky130_fd_sc_hd__clkbuf_1 _12995_ (.A(_06552_),
    .X(_00939_));
 sky130_fd_sc_hd__mux2_1 _12996_ (.A0(_05263_),
    .A1(\regs[20][12] ),
    .S(_06550_),
    .X(_06553_));
 sky130_fd_sc_hd__clkbuf_1 _12997_ (.A(_06553_),
    .X(_00940_));
 sky130_fd_sc_hd__mux2_1 _12998_ (.A0(_05296_),
    .A1(\regs[20][13] ),
    .S(_06550_),
    .X(_06554_));
 sky130_fd_sc_hd__clkbuf_1 _12999_ (.A(_06554_),
    .X(_00941_));
 sky130_fd_sc_hd__mux2_1 _13000_ (.A0(_05329_),
    .A1(\regs[20][14] ),
    .S(_06550_),
    .X(_06555_));
 sky130_fd_sc_hd__clkbuf_1 _13001_ (.A(_06555_),
    .X(_00942_));
 sky130_fd_sc_hd__mux2_1 _13002_ (.A0(_05359_),
    .A1(\regs[20][15] ),
    .S(_06550_),
    .X(_06556_));
 sky130_fd_sc_hd__clkbuf_1 _13003_ (.A(_06556_),
    .X(_00943_));
 sky130_fd_sc_hd__mux2_1 _13004_ (.A0(_05400_),
    .A1(\regs[20][16] ),
    .S(_06550_),
    .X(_06557_));
 sky130_fd_sc_hd__clkbuf_1 _13005_ (.A(_06557_),
    .X(_00944_));
 sky130_fd_sc_hd__mux2_1 _13006_ (.A0(_05424_),
    .A1(\regs[20][17] ),
    .S(_06550_),
    .X(_06558_));
 sky130_fd_sc_hd__clkbuf_1 _13007_ (.A(_06558_),
    .X(_00945_));
 sky130_fd_sc_hd__mux2_1 _13008_ (.A0(_05452_),
    .A1(\regs[20][18] ),
    .S(_06550_),
    .X(_06559_));
 sky130_fd_sc_hd__clkbuf_1 _13009_ (.A(_06559_),
    .X(_00946_));
 sky130_fd_sc_hd__mux2_1 _13010_ (.A0(_05477_),
    .A1(\regs[20][19] ),
    .S(_06550_),
    .X(_06560_));
 sky130_fd_sc_hd__clkbuf_1 _13011_ (.A(_06560_),
    .X(_00947_));
 sky130_fd_sc_hd__buf_6 _13012_ (.A(_06538_),
    .X(_06561_));
 sky130_fd_sc_hd__mux2_1 _13013_ (.A0(_05514_),
    .A1(\regs[20][20] ),
    .S(_06561_),
    .X(_06562_));
 sky130_fd_sc_hd__clkbuf_1 _13014_ (.A(_06562_),
    .X(_00948_));
 sky130_fd_sc_hd__mux2_1 _13015_ (.A0(_05541_),
    .A1(\regs[20][21] ),
    .S(_06561_),
    .X(_06563_));
 sky130_fd_sc_hd__clkbuf_1 _13016_ (.A(_06563_),
    .X(_00949_));
 sky130_fd_sc_hd__mux2_1 _13017_ (.A0(_05570_),
    .A1(\regs[20][22] ),
    .S(_06561_),
    .X(_06564_));
 sky130_fd_sc_hd__clkbuf_1 _13018_ (.A(_06564_),
    .X(_00950_));
 sky130_fd_sc_hd__mux2_1 _13019_ (.A0(_05600_),
    .A1(\regs[20][23] ),
    .S(_06561_),
    .X(_06565_));
 sky130_fd_sc_hd__clkbuf_1 _13020_ (.A(_06565_),
    .X(_00951_));
 sky130_fd_sc_hd__mux2_1 _13021_ (.A0(_05636_),
    .A1(\regs[20][24] ),
    .S(_06561_),
    .X(_06566_));
 sky130_fd_sc_hd__clkbuf_1 _13022_ (.A(_06566_),
    .X(_00952_));
 sky130_fd_sc_hd__mux2_1 _13023_ (.A0(_05660_),
    .A1(\regs[20][25] ),
    .S(_06561_),
    .X(_06567_));
 sky130_fd_sc_hd__clkbuf_1 _13024_ (.A(_06567_),
    .X(_00953_));
 sky130_fd_sc_hd__mux2_1 _13025_ (.A0(_05684_),
    .A1(\regs[20][26] ),
    .S(_06561_),
    .X(_06568_));
 sky130_fd_sc_hd__clkbuf_1 _13026_ (.A(_06568_),
    .X(_00954_));
 sky130_fd_sc_hd__mux2_1 _13027_ (.A0(_05708_),
    .A1(\regs[20][27] ),
    .S(_06561_),
    .X(_06569_));
 sky130_fd_sc_hd__clkbuf_1 _13028_ (.A(_06569_),
    .X(_00955_));
 sky130_fd_sc_hd__mux2_1 _13029_ (.A0(_05735_),
    .A1(\regs[20][28] ),
    .S(_06561_),
    .X(_06570_));
 sky130_fd_sc_hd__clkbuf_1 _13030_ (.A(_06570_),
    .X(_00956_));
 sky130_fd_sc_hd__mux2_1 _13031_ (.A0(_05763_),
    .A1(\regs[20][29] ),
    .S(_06561_),
    .X(_06571_));
 sky130_fd_sc_hd__clkbuf_1 _13032_ (.A(_06571_),
    .X(_00957_));
 sky130_fd_sc_hd__mux2_1 _13033_ (.A0(_05787_),
    .A1(\regs[20][30] ),
    .S(_06538_),
    .X(_06572_));
 sky130_fd_sc_hd__clkbuf_1 _13034_ (.A(_06572_),
    .X(_00958_));
 sky130_fd_sc_hd__mux2_1 _13035_ (.A0(_05811_),
    .A1(\regs[20][31] ),
    .S(_06538_),
    .X(_06573_));
 sky130_fd_sc_hd__clkbuf_1 _13036_ (.A(_06573_),
    .X(_00959_));
 sky130_fd_sc_hd__nor2_4 _13037_ (.A(_06072_),
    .B(_06537_),
    .Y(_06574_));
 sky130_fd_sc_hd__buf_6 _13038_ (.A(_06574_),
    .X(_06575_));
 sky130_fd_sc_hd__mux2_1 _13039_ (.A0(\regs[21][0] ),
    .A1(_06291_),
    .S(_06575_),
    .X(_06576_));
 sky130_fd_sc_hd__clkbuf_1 _13040_ (.A(_06576_),
    .X(_00960_));
 sky130_fd_sc_hd__mux2_1 _13041_ (.A0(\regs[21][1] ),
    .A1(_06295_),
    .S(_06575_),
    .X(_06577_));
 sky130_fd_sc_hd__clkbuf_1 _13042_ (.A(_06577_),
    .X(_00961_));
 sky130_fd_sc_hd__mux2_1 _13043_ (.A0(\regs[21][2] ),
    .A1(_06297_),
    .S(_06575_),
    .X(_06578_));
 sky130_fd_sc_hd__clkbuf_1 _13044_ (.A(_06578_),
    .X(_00962_));
 sky130_fd_sc_hd__mux2_1 _13045_ (.A0(\regs[21][3] ),
    .A1(_06299_),
    .S(_06575_),
    .X(_06579_));
 sky130_fd_sc_hd__clkbuf_1 _13046_ (.A(_06579_),
    .X(_00963_));
 sky130_fd_sc_hd__mux2_1 _13047_ (.A0(\regs[21][4] ),
    .A1(_06301_),
    .S(_06575_),
    .X(_06580_));
 sky130_fd_sc_hd__clkbuf_1 _13048_ (.A(_06580_),
    .X(_00964_));
 sky130_fd_sc_hd__mux2_1 _13049_ (.A0(\regs[21][5] ),
    .A1(_06303_),
    .S(_06575_),
    .X(_06581_));
 sky130_fd_sc_hd__clkbuf_1 _13050_ (.A(_06581_),
    .X(_00965_));
 sky130_fd_sc_hd__mux2_1 _13051_ (.A0(\regs[21][6] ),
    .A1(_06305_),
    .S(_06575_),
    .X(_06582_));
 sky130_fd_sc_hd__clkbuf_1 _13052_ (.A(_06582_),
    .X(_00966_));
 sky130_fd_sc_hd__mux2_1 _13053_ (.A0(\regs[21][7] ),
    .A1(_06307_),
    .S(_06575_),
    .X(_06583_));
 sky130_fd_sc_hd__clkbuf_1 _13054_ (.A(_06583_),
    .X(_00967_));
 sky130_fd_sc_hd__mux2_1 _13055_ (.A0(\regs[21][8] ),
    .A1(_06309_),
    .S(_06575_),
    .X(_06584_));
 sky130_fd_sc_hd__clkbuf_1 _13056_ (.A(_06584_),
    .X(_00968_));
 sky130_fd_sc_hd__mux2_1 _13057_ (.A0(\regs[21][9] ),
    .A1(_06311_),
    .S(_06575_),
    .X(_06585_));
 sky130_fd_sc_hd__clkbuf_1 _13058_ (.A(_06585_),
    .X(_00969_));
 sky130_fd_sc_hd__buf_6 _13059_ (.A(_06574_),
    .X(_06586_));
 sky130_fd_sc_hd__mux2_1 _13060_ (.A0(\regs[21][10] ),
    .A1(_06313_),
    .S(_06586_),
    .X(_06587_));
 sky130_fd_sc_hd__clkbuf_1 _13061_ (.A(_06587_),
    .X(_00970_));
 sky130_fd_sc_hd__mux2_1 _13062_ (.A0(\regs[21][11] ),
    .A1(_06316_),
    .S(_06586_),
    .X(_06588_));
 sky130_fd_sc_hd__clkbuf_1 _13063_ (.A(_06588_),
    .X(_00971_));
 sky130_fd_sc_hd__mux2_1 _13064_ (.A0(\regs[21][12] ),
    .A1(_06318_),
    .S(_06586_),
    .X(_06589_));
 sky130_fd_sc_hd__clkbuf_1 _13065_ (.A(_06589_),
    .X(_00972_));
 sky130_fd_sc_hd__mux2_1 _13066_ (.A0(\regs[21][13] ),
    .A1(_06320_),
    .S(_06586_),
    .X(_06590_));
 sky130_fd_sc_hd__clkbuf_1 _13067_ (.A(_06590_),
    .X(_00973_));
 sky130_fd_sc_hd__mux2_1 _13068_ (.A0(\regs[21][14] ),
    .A1(_06322_),
    .S(_06586_),
    .X(_06591_));
 sky130_fd_sc_hd__clkbuf_1 _13069_ (.A(_06591_),
    .X(_00974_));
 sky130_fd_sc_hd__mux2_1 _13070_ (.A0(\regs[21][15] ),
    .A1(_06324_),
    .S(_06586_),
    .X(_06592_));
 sky130_fd_sc_hd__clkbuf_1 _13071_ (.A(_06592_),
    .X(_00975_));
 sky130_fd_sc_hd__mux2_1 _13072_ (.A0(\regs[21][16] ),
    .A1(_06326_),
    .S(_06586_),
    .X(_06593_));
 sky130_fd_sc_hd__clkbuf_1 _13073_ (.A(_06593_),
    .X(_00976_));
 sky130_fd_sc_hd__mux2_1 _13074_ (.A0(\regs[21][17] ),
    .A1(_06328_),
    .S(_06586_),
    .X(_06594_));
 sky130_fd_sc_hd__clkbuf_1 _13075_ (.A(_06594_),
    .X(_00977_));
 sky130_fd_sc_hd__mux2_1 _13076_ (.A0(\regs[21][18] ),
    .A1(_06330_),
    .S(_06586_),
    .X(_06595_));
 sky130_fd_sc_hd__clkbuf_1 _13077_ (.A(_06595_),
    .X(_00978_));
 sky130_fd_sc_hd__mux2_1 _13078_ (.A0(\regs[21][19] ),
    .A1(_06332_),
    .S(_06586_),
    .X(_06596_));
 sky130_fd_sc_hd__clkbuf_1 _13079_ (.A(_06596_),
    .X(_00979_));
 sky130_fd_sc_hd__buf_4 _13080_ (.A(_06574_),
    .X(_06597_));
 sky130_fd_sc_hd__mux2_1 _13081_ (.A0(\regs[21][20] ),
    .A1(_06334_),
    .S(_06597_),
    .X(_06598_));
 sky130_fd_sc_hd__clkbuf_1 _13082_ (.A(_06598_),
    .X(_00980_));
 sky130_fd_sc_hd__mux2_1 _13083_ (.A0(\regs[21][21] ),
    .A1(_06337_),
    .S(_06597_),
    .X(_06599_));
 sky130_fd_sc_hd__clkbuf_1 _13084_ (.A(_06599_),
    .X(_00981_));
 sky130_fd_sc_hd__mux2_1 _13085_ (.A0(\regs[21][22] ),
    .A1(_06339_),
    .S(_06597_),
    .X(_06600_));
 sky130_fd_sc_hd__clkbuf_1 _13086_ (.A(_06600_),
    .X(_00982_));
 sky130_fd_sc_hd__mux2_1 _13087_ (.A0(\regs[21][23] ),
    .A1(_06341_),
    .S(_06597_),
    .X(_06601_));
 sky130_fd_sc_hd__clkbuf_1 _13088_ (.A(_06601_),
    .X(_00983_));
 sky130_fd_sc_hd__mux2_1 _13089_ (.A0(\regs[21][24] ),
    .A1(_06343_),
    .S(_06597_),
    .X(_06602_));
 sky130_fd_sc_hd__clkbuf_1 _13090_ (.A(_06602_),
    .X(_00984_));
 sky130_fd_sc_hd__mux2_1 _13091_ (.A0(\regs[21][25] ),
    .A1(_06345_),
    .S(_06597_),
    .X(_06603_));
 sky130_fd_sc_hd__clkbuf_1 _13092_ (.A(_06603_),
    .X(_00985_));
 sky130_fd_sc_hd__mux2_1 _13093_ (.A0(\regs[21][26] ),
    .A1(_06347_),
    .S(_06597_),
    .X(_06604_));
 sky130_fd_sc_hd__clkbuf_1 _13094_ (.A(_06604_),
    .X(_00986_));
 sky130_fd_sc_hd__mux2_1 _13095_ (.A0(\regs[21][27] ),
    .A1(_06349_),
    .S(_06597_),
    .X(_06605_));
 sky130_fd_sc_hd__clkbuf_1 _13096_ (.A(_06605_),
    .X(_00987_));
 sky130_fd_sc_hd__mux2_1 _13097_ (.A0(\regs[21][28] ),
    .A1(_06351_),
    .S(_06597_),
    .X(_06606_));
 sky130_fd_sc_hd__clkbuf_1 _13098_ (.A(_06606_),
    .X(_00988_));
 sky130_fd_sc_hd__mux2_1 _13099_ (.A0(\regs[21][29] ),
    .A1(_06353_),
    .S(_06597_),
    .X(_06607_));
 sky130_fd_sc_hd__clkbuf_1 _13100_ (.A(_06607_),
    .X(_00989_));
 sky130_fd_sc_hd__mux2_1 _13101_ (.A0(\regs[21][30] ),
    .A1(_06355_),
    .S(_06574_),
    .X(_06608_));
 sky130_fd_sc_hd__clkbuf_1 _13102_ (.A(_06608_),
    .X(_00990_));
 sky130_fd_sc_hd__mux2_1 _13103_ (.A0(\regs[21][31] ),
    .A1(_06357_),
    .S(_06574_),
    .X(_06609_));
 sky130_fd_sc_hd__clkbuf_1 _13104_ (.A(_06609_),
    .X(_00991_));
 sky130_fd_sc_hd__nor2_4 _13105_ (.A(_05883_),
    .B(_06537_),
    .Y(_06610_));
 sky130_fd_sc_hd__buf_6 _13106_ (.A(_06610_),
    .X(_06611_));
 sky130_fd_sc_hd__mux2_1 _13107_ (.A0(\regs[22][0] ),
    .A1(_06291_),
    .S(_06611_),
    .X(_06612_));
 sky130_fd_sc_hd__clkbuf_1 _13108_ (.A(_06612_),
    .X(_00992_));
 sky130_fd_sc_hd__mux2_1 _13109_ (.A0(\regs[22][1] ),
    .A1(_06295_),
    .S(_06611_),
    .X(_06613_));
 sky130_fd_sc_hd__clkbuf_1 _13110_ (.A(_06613_),
    .X(_00993_));
 sky130_fd_sc_hd__mux2_1 _13111_ (.A0(\regs[22][2] ),
    .A1(_06297_),
    .S(_06611_),
    .X(_06614_));
 sky130_fd_sc_hd__clkbuf_1 _13112_ (.A(_06614_),
    .X(_00994_));
 sky130_fd_sc_hd__mux2_1 _13113_ (.A0(\regs[22][3] ),
    .A1(_06299_),
    .S(_06611_),
    .X(_06615_));
 sky130_fd_sc_hd__clkbuf_1 _13114_ (.A(_06615_),
    .X(_00995_));
 sky130_fd_sc_hd__mux2_1 _13115_ (.A0(\regs[22][4] ),
    .A1(_06301_),
    .S(_06611_),
    .X(_06616_));
 sky130_fd_sc_hd__clkbuf_1 _13116_ (.A(_06616_),
    .X(_00996_));
 sky130_fd_sc_hd__mux2_1 _13117_ (.A0(\regs[22][5] ),
    .A1(_06303_),
    .S(_06611_),
    .X(_06617_));
 sky130_fd_sc_hd__clkbuf_1 _13118_ (.A(_06617_),
    .X(_00997_));
 sky130_fd_sc_hd__mux2_1 _13119_ (.A0(\regs[22][6] ),
    .A1(_06305_),
    .S(_06611_),
    .X(_06618_));
 sky130_fd_sc_hd__clkbuf_1 _13120_ (.A(_06618_),
    .X(_00998_));
 sky130_fd_sc_hd__mux2_1 _13121_ (.A0(\regs[22][7] ),
    .A1(_06307_),
    .S(_06611_),
    .X(_06619_));
 sky130_fd_sc_hd__clkbuf_1 _13122_ (.A(_06619_),
    .X(_00999_));
 sky130_fd_sc_hd__mux2_1 _13123_ (.A0(\regs[22][8] ),
    .A1(_06309_),
    .S(_06611_),
    .X(_06620_));
 sky130_fd_sc_hd__clkbuf_1 _13124_ (.A(_06620_),
    .X(_01000_));
 sky130_fd_sc_hd__mux2_1 _13125_ (.A0(\regs[22][9] ),
    .A1(_06311_),
    .S(_06611_),
    .X(_06621_));
 sky130_fd_sc_hd__clkbuf_1 _13126_ (.A(_06621_),
    .X(_01001_));
 sky130_fd_sc_hd__buf_6 _13127_ (.A(_06610_),
    .X(_06622_));
 sky130_fd_sc_hd__mux2_1 _13128_ (.A0(\regs[22][10] ),
    .A1(_06313_),
    .S(_06622_),
    .X(_06623_));
 sky130_fd_sc_hd__clkbuf_1 _13129_ (.A(_06623_),
    .X(_01002_));
 sky130_fd_sc_hd__mux2_1 _13130_ (.A0(\regs[22][11] ),
    .A1(_06316_),
    .S(_06622_),
    .X(_06624_));
 sky130_fd_sc_hd__clkbuf_1 _13131_ (.A(_06624_),
    .X(_01003_));
 sky130_fd_sc_hd__mux2_1 _13132_ (.A0(\regs[22][12] ),
    .A1(_06318_),
    .S(_06622_),
    .X(_06625_));
 sky130_fd_sc_hd__clkbuf_1 _13133_ (.A(_06625_),
    .X(_01004_));
 sky130_fd_sc_hd__mux2_1 _13134_ (.A0(\regs[22][13] ),
    .A1(_06320_),
    .S(_06622_),
    .X(_06626_));
 sky130_fd_sc_hd__clkbuf_1 _13135_ (.A(_06626_),
    .X(_01005_));
 sky130_fd_sc_hd__mux2_1 _13136_ (.A0(\regs[22][14] ),
    .A1(_06322_),
    .S(_06622_),
    .X(_06627_));
 sky130_fd_sc_hd__clkbuf_1 _13137_ (.A(_06627_),
    .X(_01006_));
 sky130_fd_sc_hd__mux2_1 _13138_ (.A0(\regs[22][15] ),
    .A1(_06324_),
    .S(_06622_),
    .X(_06628_));
 sky130_fd_sc_hd__clkbuf_1 _13139_ (.A(_06628_),
    .X(_01007_));
 sky130_fd_sc_hd__mux2_1 _13140_ (.A0(\regs[22][16] ),
    .A1(_06326_),
    .S(_06622_),
    .X(_06629_));
 sky130_fd_sc_hd__clkbuf_1 _13141_ (.A(_06629_),
    .X(_01008_));
 sky130_fd_sc_hd__mux2_1 _13142_ (.A0(\regs[22][17] ),
    .A1(_06328_),
    .S(_06622_),
    .X(_06630_));
 sky130_fd_sc_hd__clkbuf_1 _13143_ (.A(_06630_),
    .X(_01009_));
 sky130_fd_sc_hd__mux2_1 _13144_ (.A0(\regs[22][18] ),
    .A1(_06330_),
    .S(_06622_),
    .X(_06631_));
 sky130_fd_sc_hd__clkbuf_1 _13145_ (.A(_06631_),
    .X(_01010_));
 sky130_fd_sc_hd__mux2_1 _13146_ (.A0(\regs[22][19] ),
    .A1(_06332_),
    .S(_06622_),
    .X(_06632_));
 sky130_fd_sc_hd__clkbuf_1 _13147_ (.A(_06632_),
    .X(_01011_));
 sky130_fd_sc_hd__clkbuf_8 _13148_ (.A(_06610_),
    .X(_06633_));
 sky130_fd_sc_hd__mux2_1 _13149_ (.A0(\regs[22][20] ),
    .A1(_06334_),
    .S(_06633_),
    .X(_06634_));
 sky130_fd_sc_hd__clkbuf_1 _13150_ (.A(_06634_),
    .X(_01012_));
 sky130_fd_sc_hd__mux2_1 _13151_ (.A0(\regs[22][21] ),
    .A1(_06337_),
    .S(_06633_),
    .X(_06635_));
 sky130_fd_sc_hd__clkbuf_1 _13152_ (.A(_06635_),
    .X(_01013_));
 sky130_fd_sc_hd__mux2_1 _13153_ (.A0(\regs[22][22] ),
    .A1(_06339_),
    .S(_06633_),
    .X(_06636_));
 sky130_fd_sc_hd__clkbuf_1 _13154_ (.A(_06636_),
    .X(_01014_));
 sky130_fd_sc_hd__mux2_1 _13155_ (.A0(\regs[22][23] ),
    .A1(_06341_),
    .S(_06633_),
    .X(_06637_));
 sky130_fd_sc_hd__clkbuf_1 _13156_ (.A(_06637_),
    .X(_01015_));
 sky130_fd_sc_hd__mux2_1 _13157_ (.A0(\regs[22][24] ),
    .A1(_06343_),
    .S(_06633_),
    .X(_06638_));
 sky130_fd_sc_hd__clkbuf_1 _13158_ (.A(_06638_),
    .X(_01016_));
 sky130_fd_sc_hd__mux2_1 _13159_ (.A0(\regs[22][25] ),
    .A1(_06345_),
    .S(_06633_),
    .X(_06639_));
 sky130_fd_sc_hd__clkbuf_1 _13160_ (.A(_06639_),
    .X(_01017_));
 sky130_fd_sc_hd__mux2_1 _13161_ (.A0(\regs[22][26] ),
    .A1(_06347_),
    .S(_06633_),
    .X(_06640_));
 sky130_fd_sc_hd__clkbuf_1 _13162_ (.A(_06640_),
    .X(_01018_));
 sky130_fd_sc_hd__mux2_1 _13163_ (.A0(\regs[22][27] ),
    .A1(_06349_),
    .S(_06633_),
    .X(_06641_));
 sky130_fd_sc_hd__clkbuf_1 _13164_ (.A(_06641_),
    .X(_01019_));
 sky130_fd_sc_hd__mux2_1 _13165_ (.A0(\regs[22][28] ),
    .A1(_06351_),
    .S(_06633_),
    .X(_06642_));
 sky130_fd_sc_hd__clkbuf_1 _13166_ (.A(_06642_),
    .X(_01020_));
 sky130_fd_sc_hd__mux2_1 _13167_ (.A0(\regs[22][29] ),
    .A1(_06353_),
    .S(_06633_),
    .X(_06643_));
 sky130_fd_sc_hd__clkbuf_1 _13168_ (.A(_06643_),
    .X(_01021_));
 sky130_fd_sc_hd__mux2_1 _13169_ (.A0(\regs[22][30] ),
    .A1(_06355_),
    .S(_06610_),
    .X(_06644_));
 sky130_fd_sc_hd__clkbuf_1 _13170_ (.A(_06644_),
    .X(_01022_));
 sky130_fd_sc_hd__mux2_1 _13171_ (.A0(\regs[22][31] ),
    .A1(_06357_),
    .S(_06610_),
    .X(_06645_));
 sky130_fd_sc_hd__clkbuf_1 _13172_ (.A(_06645_),
    .X(_01023_));
 sky130_fd_sc_hd__nor2_4 _13173_ (.A(_05958_),
    .B(_06537_),
    .Y(_06646_));
 sky130_fd_sc_hd__buf_6 _13174_ (.A(_06646_),
    .X(_06647_));
 sky130_fd_sc_hd__mux2_1 _13175_ (.A0(\regs[23][0] ),
    .A1(_06291_),
    .S(_06647_),
    .X(_06648_));
 sky130_fd_sc_hd__clkbuf_1 _13176_ (.A(_06648_),
    .X(_01024_));
 sky130_fd_sc_hd__mux2_1 _13177_ (.A0(\regs[23][1] ),
    .A1(_06295_),
    .S(_06647_),
    .X(_06649_));
 sky130_fd_sc_hd__clkbuf_1 _13178_ (.A(_06649_),
    .X(_01025_));
 sky130_fd_sc_hd__mux2_1 _13179_ (.A0(\regs[23][2] ),
    .A1(_06297_),
    .S(_06647_),
    .X(_06650_));
 sky130_fd_sc_hd__clkbuf_1 _13180_ (.A(_06650_),
    .X(_01026_));
 sky130_fd_sc_hd__mux2_1 _13181_ (.A0(\regs[23][3] ),
    .A1(_06299_),
    .S(_06647_),
    .X(_06651_));
 sky130_fd_sc_hd__clkbuf_1 _13182_ (.A(_06651_),
    .X(_01027_));
 sky130_fd_sc_hd__mux2_1 _13183_ (.A0(\regs[23][4] ),
    .A1(_06301_),
    .S(_06647_),
    .X(_06652_));
 sky130_fd_sc_hd__clkbuf_1 _13184_ (.A(_06652_),
    .X(_01028_));
 sky130_fd_sc_hd__mux2_1 _13185_ (.A0(\regs[23][5] ),
    .A1(_06303_),
    .S(_06647_),
    .X(_06653_));
 sky130_fd_sc_hd__clkbuf_1 _13186_ (.A(_06653_),
    .X(_01029_));
 sky130_fd_sc_hd__mux2_1 _13187_ (.A0(\regs[23][6] ),
    .A1(_06305_),
    .S(_06647_),
    .X(_06654_));
 sky130_fd_sc_hd__clkbuf_1 _13188_ (.A(_06654_),
    .X(_01030_));
 sky130_fd_sc_hd__mux2_1 _13189_ (.A0(\regs[23][7] ),
    .A1(_06307_),
    .S(_06647_),
    .X(_06655_));
 sky130_fd_sc_hd__clkbuf_1 _13190_ (.A(_06655_),
    .X(_01031_));
 sky130_fd_sc_hd__mux2_1 _13191_ (.A0(\regs[23][8] ),
    .A1(_06309_),
    .S(_06647_),
    .X(_06656_));
 sky130_fd_sc_hd__clkbuf_1 _13192_ (.A(_06656_),
    .X(_01032_));
 sky130_fd_sc_hd__mux2_1 _13193_ (.A0(\regs[23][9] ),
    .A1(_06311_),
    .S(_06647_),
    .X(_06657_));
 sky130_fd_sc_hd__clkbuf_1 _13194_ (.A(_06657_),
    .X(_01033_));
 sky130_fd_sc_hd__clkbuf_8 _13195_ (.A(_06646_),
    .X(_06658_));
 sky130_fd_sc_hd__mux2_1 _13196_ (.A0(\regs[23][10] ),
    .A1(_06313_),
    .S(_06658_),
    .X(_06659_));
 sky130_fd_sc_hd__clkbuf_1 _13197_ (.A(_06659_),
    .X(_01034_));
 sky130_fd_sc_hd__mux2_1 _13198_ (.A0(\regs[23][11] ),
    .A1(_06316_),
    .S(_06658_),
    .X(_06660_));
 sky130_fd_sc_hd__clkbuf_1 _13199_ (.A(_06660_),
    .X(_01035_));
 sky130_fd_sc_hd__mux2_1 _13200_ (.A0(\regs[23][12] ),
    .A1(_06318_),
    .S(_06658_),
    .X(_06661_));
 sky130_fd_sc_hd__clkbuf_1 _13201_ (.A(_06661_),
    .X(_01036_));
 sky130_fd_sc_hd__mux2_1 _13202_ (.A0(\regs[23][13] ),
    .A1(_06320_),
    .S(_06658_),
    .X(_06662_));
 sky130_fd_sc_hd__clkbuf_1 _13203_ (.A(_06662_),
    .X(_01037_));
 sky130_fd_sc_hd__mux2_1 _13204_ (.A0(\regs[23][14] ),
    .A1(_06322_),
    .S(_06658_),
    .X(_06663_));
 sky130_fd_sc_hd__clkbuf_1 _13205_ (.A(_06663_),
    .X(_01038_));
 sky130_fd_sc_hd__mux2_1 _13206_ (.A0(\regs[23][15] ),
    .A1(_06324_),
    .S(_06658_),
    .X(_06664_));
 sky130_fd_sc_hd__clkbuf_1 _13207_ (.A(_06664_),
    .X(_01039_));
 sky130_fd_sc_hd__mux2_1 _13208_ (.A0(\regs[23][16] ),
    .A1(_06326_),
    .S(_06658_),
    .X(_06665_));
 sky130_fd_sc_hd__clkbuf_1 _13209_ (.A(_06665_),
    .X(_01040_));
 sky130_fd_sc_hd__mux2_1 _13210_ (.A0(\regs[23][17] ),
    .A1(_06328_),
    .S(_06658_),
    .X(_06666_));
 sky130_fd_sc_hd__clkbuf_1 _13211_ (.A(_06666_),
    .X(_01041_));
 sky130_fd_sc_hd__mux2_1 _13212_ (.A0(\regs[23][18] ),
    .A1(_06330_),
    .S(_06658_),
    .X(_06667_));
 sky130_fd_sc_hd__clkbuf_1 _13213_ (.A(_06667_),
    .X(_01042_));
 sky130_fd_sc_hd__mux2_1 _13214_ (.A0(\regs[23][19] ),
    .A1(_06332_),
    .S(_06658_),
    .X(_06668_));
 sky130_fd_sc_hd__clkbuf_1 _13215_ (.A(_06668_),
    .X(_01043_));
 sky130_fd_sc_hd__clkbuf_8 _13216_ (.A(_06646_),
    .X(_06669_));
 sky130_fd_sc_hd__mux2_1 _13217_ (.A0(\regs[23][20] ),
    .A1(_06334_),
    .S(_06669_),
    .X(_06670_));
 sky130_fd_sc_hd__clkbuf_1 _13218_ (.A(_06670_),
    .X(_01044_));
 sky130_fd_sc_hd__mux2_1 _13219_ (.A0(\regs[23][21] ),
    .A1(_06337_),
    .S(_06669_),
    .X(_06671_));
 sky130_fd_sc_hd__clkbuf_1 _13220_ (.A(_06671_),
    .X(_01045_));
 sky130_fd_sc_hd__mux2_1 _13221_ (.A0(\regs[23][22] ),
    .A1(_06339_),
    .S(_06669_),
    .X(_06672_));
 sky130_fd_sc_hd__clkbuf_1 _13222_ (.A(_06672_),
    .X(_01046_));
 sky130_fd_sc_hd__mux2_1 _13223_ (.A0(\regs[23][23] ),
    .A1(_06341_),
    .S(_06669_),
    .X(_06673_));
 sky130_fd_sc_hd__clkbuf_1 _13224_ (.A(_06673_),
    .X(_01047_));
 sky130_fd_sc_hd__mux2_1 _13225_ (.A0(\regs[23][24] ),
    .A1(_06343_),
    .S(_06669_),
    .X(_06674_));
 sky130_fd_sc_hd__clkbuf_1 _13226_ (.A(_06674_),
    .X(_01048_));
 sky130_fd_sc_hd__mux2_1 _13227_ (.A0(\regs[23][25] ),
    .A1(_06345_),
    .S(_06669_),
    .X(_06675_));
 sky130_fd_sc_hd__clkbuf_1 _13228_ (.A(_06675_),
    .X(_01049_));
 sky130_fd_sc_hd__mux2_1 _13229_ (.A0(\regs[23][26] ),
    .A1(_06347_),
    .S(_06669_),
    .X(_06676_));
 sky130_fd_sc_hd__clkbuf_1 _13230_ (.A(_06676_),
    .X(_01050_));
 sky130_fd_sc_hd__mux2_1 _13231_ (.A0(\regs[23][27] ),
    .A1(_06349_),
    .S(_06669_),
    .X(_06677_));
 sky130_fd_sc_hd__clkbuf_1 _13232_ (.A(_06677_),
    .X(_01051_));
 sky130_fd_sc_hd__mux2_1 _13233_ (.A0(\regs[23][28] ),
    .A1(_06351_),
    .S(_06669_),
    .X(_06678_));
 sky130_fd_sc_hd__clkbuf_1 _13234_ (.A(_06678_),
    .X(_01052_));
 sky130_fd_sc_hd__mux2_1 _13235_ (.A0(\regs[23][29] ),
    .A1(_06353_),
    .S(_06669_),
    .X(_06679_));
 sky130_fd_sc_hd__clkbuf_1 _13236_ (.A(_06679_),
    .X(_01053_));
 sky130_fd_sc_hd__mux2_1 _13237_ (.A0(\regs[23][30] ),
    .A1(_06355_),
    .S(_06646_),
    .X(_06680_));
 sky130_fd_sc_hd__clkbuf_1 _13238_ (.A(_06680_),
    .X(_01054_));
 sky130_fd_sc_hd__mux2_1 _13239_ (.A0(\regs[23][31] ),
    .A1(_06357_),
    .S(_06646_),
    .X(_06681_));
 sky130_fd_sc_hd__clkbuf_1 _13240_ (.A(_06681_),
    .X(_01055_));
 sky130_fd_sc_hd__and4b_2 _13241_ (.A_N(_02241_),
    .B(_04765_),
    .C(_02313_),
    .D(_02315_),
    .X(_06682_));
 sky130_fd_sc_hd__nand2_2 _13242_ (.A(_06031_),
    .B(_06682_),
    .Y(_06683_));
 sky130_fd_sc_hd__buf_4 _13243_ (.A(_06683_),
    .X(_06684_));
 sky130_fd_sc_hd__mux2_1 _13244_ (.A0(_04762_),
    .A1(\regs[24][0] ),
    .S(_06684_),
    .X(_06685_));
 sky130_fd_sc_hd__clkbuf_1 _13245_ (.A(_06685_),
    .X(_01056_));
 sky130_fd_sc_hd__mux2_1 _13246_ (.A0(_04818_),
    .A1(\regs[24][1] ),
    .S(_06684_),
    .X(_06686_));
 sky130_fd_sc_hd__clkbuf_1 _13247_ (.A(_06686_),
    .X(_01057_));
 sky130_fd_sc_hd__mux2_1 _13248_ (.A0(_04858_),
    .A1(\regs[24][2] ),
    .S(_06684_),
    .X(_06687_));
 sky130_fd_sc_hd__clkbuf_1 _13249_ (.A(_06687_),
    .X(_01058_));
 sky130_fd_sc_hd__mux2_1 _13250_ (.A0(_04904_),
    .A1(\regs[24][3] ),
    .S(_06684_),
    .X(_06688_));
 sky130_fd_sc_hd__clkbuf_1 _13251_ (.A(_06688_),
    .X(_01059_));
 sky130_fd_sc_hd__mux2_1 _13252_ (.A0(_04952_),
    .A1(\regs[24][4] ),
    .S(_06684_),
    .X(_06689_));
 sky130_fd_sc_hd__clkbuf_1 _13253_ (.A(_06689_),
    .X(_01060_));
 sky130_fd_sc_hd__mux2_1 _13254_ (.A0(_04992_),
    .A1(\regs[24][5] ),
    .S(_06684_),
    .X(_06690_));
 sky130_fd_sc_hd__clkbuf_1 _13255_ (.A(_06690_),
    .X(_01061_));
 sky130_fd_sc_hd__mux2_1 _13256_ (.A0(_05030_),
    .A1(\regs[24][6] ),
    .S(_06684_),
    .X(_06691_));
 sky130_fd_sc_hd__clkbuf_1 _13257_ (.A(_06691_),
    .X(_01062_));
 sky130_fd_sc_hd__mux2_1 _13258_ (.A0(_05080_),
    .A1(\regs[24][7] ),
    .S(_06684_),
    .X(_06692_));
 sky130_fd_sc_hd__clkbuf_1 _13259_ (.A(_06692_),
    .X(_01063_));
 sky130_fd_sc_hd__mux2_1 _13260_ (.A0(_05121_),
    .A1(\regs[24][8] ),
    .S(_06684_),
    .X(_06693_));
 sky130_fd_sc_hd__clkbuf_1 _13261_ (.A(_06693_),
    .X(_01064_));
 sky130_fd_sc_hd__mux2_1 _13262_ (.A0(_05157_),
    .A1(\regs[24][9] ),
    .S(_06684_),
    .X(_06694_));
 sky130_fd_sc_hd__clkbuf_1 _13263_ (.A(_06694_),
    .X(_01065_));
 sky130_fd_sc_hd__buf_6 _13264_ (.A(_06683_),
    .X(_06695_));
 sky130_fd_sc_hd__mux2_1 _13265_ (.A0(_05187_),
    .A1(\regs[24][10] ),
    .S(_06695_),
    .X(_06696_));
 sky130_fd_sc_hd__clkbuf_1 _13266_ (.A(_06696_),
    .X(_01066_));
 sky130_fd_sc_hd__mux2_1 _13267_ (.A0(_05224_),
    .A1(\regs[24][11] ),
    .S(_06695_),
    .X(_06697_));
 sky130_fd_sc_hd__clkbuf_1 _13268_ (.A(_06697_),
    .X(_01067_));
 sky130_fd_sc_hd__mux2_1 _13269_ (.A0(_05263_),
    .A1(\regs[24][12] ),
    .S(_06695_),
    .X(_06698_));
 sky130_fd_sc_hd__clkbuf_1 _13270_ (.A(_06698_),
    .X(_01068_));
 sky130_fd_sc_hd__mux2_1 _13271_ (.A0(_05296_),
    .A1(\regs[24][13] ),
    .S(_06695_),
    .X(_06699_));
 sky130_fd_sc_hd__clkbuf_1 _13272_ (.A(_06699_),
    .X(_01069_));
 sky130_fd_sc_hd__mux2_1 _13273_ (.A0(_05329_),
    .A1(\regs[24][14] ),
    .S(_06695_),
    .X(_06700_));
 sky130_fd_sc_hd__clkbuf_1 _13274_ (.A(_06700_),
    .X(_01070_));
 sky130_fd_sc_hd__mux2_1 _13275_ (.A0(_05359_),
    .A1(\regs[24][15] ),
    .S(_06695_),
    .X(_06701_));
 sky130_fd_sc_hd__clkbuf_1 _13276_ (.A(_06701_),
    .X(_01071_));
 sky130_fd_sc_hd__mux2_1 _13277_ (.A0(_05400_),
    .A1(\regs[24][16] ),
    .S(_06695_),
    .X(_06702_));
 sky130_fd_sc_hd__clkbuf_1 _13278_ (.A(_06702_),
    .X(_01072_));
 sky130_fd_sc_hd__mux2_1 _13279_ (.A0(_05424_),
    .A1(\regs[24][17] ),
    .S(_06695_),
    .X(_06703_));
 sky130_fd_sc_hd__clkbuf_1 _13280_ (.A(_06703_),
    .X(_01073_));
 sky130_fd_sc_hd__mux2_1 _13281_ (.A0(_05452_),
    .A1(\regs[24][18] ),
    .S(_06695_),
    .X(_06704_));
 sky130_fd_sc_hd__clkbuf_1 _13282_ (.A(_06704_),
    .X(_01074_));
 sky130_fd_sc_hd__mux2_1 _13283_ (.A0(_05477_),
    .A1(\regs[24][19] ),
    .S(_06695_),
    .X(_06705_));
 sky130_fd_sc_hd__clkbuf_1 _13284_ (.A(_06705_),
    .X(_01075_));
 sky130_fd_sc_hd__buf_4 _13285_ (.A(_06683_),
    .X(_06706_));
 sky130_fd_sc_hd__mux2_1 _13286_ (.A0(_05514_),
    .A1(\regs[24][20] ),
    .S(_06706_),
    .X(_06707_));
 sky130_fd_sc_hd__clkbuf_1 _13287_ (.A(_06707_),
    .X(_01076_));
 sky130_fd_sc_hd__mux2_1 _13288_ (.A0(_05541_),
    .A1(\regs[24][21] ),
    .S(_06706_),
    .X(_06708_));
 sky130_fd_sc_hd__clkbuf_1 _13289_ (.A(_06708_),
    .X(_01077_));
 sky130_fd_sc_hd__mux2_1 _13290_ (.A0(_05570_),
    .A1(\regs[24][22] ),
    .S(_06706_),
    .X(_06709_));
 sky130_fd_sc_hd__clkbuf_1 _13291_ (.A(_06709_),
    .X(_01078_));
 sky130_fd_sc_hd__mux2_1 _13292_ (.A0(_05600_),
    .A1(\regs[24][23] ),
    .S(_06706_),
    .X(_06710_));
 sky130_fd_sc_hd__clkbuf_1 _13293_ (.A(_06710_),
    .X(_01079_));
 sky130_fd_sc_hd__mux2_1 _13294_ (.A0(_05636_),
    .A1(\regs[24][24] ),
    .S(_06706_),
    .X(_06711_));
 sky130_fd_sc_hd__clkbuf_1 _13295_ (.A(_06711_),
    .X(_01080_));
 sky130_fd_sc_hd__mux2_1 _13296_ (.A0(_05660_),
    .A1(\regs[24][25] ),
    .S(_06706_),
    .X(_06712_));
 sky130_fd_sc_hd__clkbuf_1 _13297_ (.A(_06712_),
    .X(_01081_));
 sky130_fd_sc_hd__mux2_1 _13298_ (.A0(_05684_),
    .A1(\regs[24][26] ),
    .S(_06706_),
    .X(_06713_));
 sky130_fd_sc_hd__clkbuf_1 _13299_ (.A(_06713_),
    .X(_01082_));
 sky130_fd_sc_hd__mux2_1 _13300_ (.A0(_05708_),
    .A1(\regs[24][27] ),
    .S(_06706_),
    .X(_06714_));
 sky130_fd_sc_hd__clkbuf_1 _13301_ (.A(_06714_),
    .X(_01083_));
 sky130_fd_sc_hd__mux2_1 _13302_ (.A0(_05735_),
    .A1(\regs[24][28] ),
    .S(_06706_),
    .X(_06715_));
 sky130_fd_sc_hd__clkbuf_1 _13303_ (.A(_06715_),
    .X(_01084_));
 sky130_fd_sc_hd__mux2_1 _13304_ (.A0(_05763_),
    .A1(\regs[24][29] ),
    .S(_06706_),
    .X(_06716_));
 sky130_fd_sc_hd__clkbuf_1 _13305_ (.A(_06716_),
    .X(_01085_));
 sky130_fd_sc_hd__mux2_1 _13306_ (.A0(_05787_),
    .A1(\regs[24][30] ),
    .S(_06683_),
    .X(_06717_));
 sky130_fd_sc_hd__clkbuf_1 _13307_ (.A(_06717_),
    .X(_01086_));
 sky130_fd_sc_hd__mux2_1 _13308_ (.A0(_05811_),
    .A1(\regs[24][31] ),
    .S(_06683_),
    .X(_06718_));
 sky130_fd_sc_hd__clkbuf_1 _13309_ (.A(_06718_),
    .X(_01087_));
 sky130_fd_sc_hd__nand2_2 _13310_ (.A(_04764_),
    .B(_06682_),
    .Y(_06719_));
 sky130_fd_sc_hd__buf_4 _13311_ (.A(_06719_),
    .X(_06720_));
 sky130_fd_sc_hd__mux2_1 _13312_ (.A0(_04762_),
    .A1(\regs[25][0] ),
    .S(_06720_),
    .X(_06721_));
 sky130_fd_sc_hd__clkbuf_1 _13313_ (.A(_06721_),
    .X(_01088_));
 sky130_fd_sc_hd__mux2_1 _13314_ (.A0(_04818_),
    .A1(\regs[25][1] ),
    .S(_06720_),
    .X(_06722_));
 sky130_fd_sc_hd__clkbuf_1 _13315_ (.A(_06722_),
    .X(_01089_));
 sky130_fd_sc_hd__mux2_1 _13316_ (.A0(_04858_),
    .A1(\regs[25][2] ),
    .S(_06720_),
    .X(_06723_));
 sky130_fd_sc_hd__clkbuf_1 _13317_ (.A(_06723_),
    .X(_01090_));
 sky130_fd_sc_hd__mux2_1 _13318_ (.A0(_04904_),
    .A1(\regs[25][3] ),
    .S(_06720_),
    .X(_06724_));
 sky130_fd_sc_hd__clkbuf_1 _13319_ (.A(_06724_),
    .X(_01091_));
 sky130_fd_sc_hd__mux2_1 _13320_ (.A0(_04952_),
    .A1(\regs[25][4] ),
    .S(_06720_),
    .X(_06725_));
 sky130_fd_sc_hd__clkbuf_1 _13321_ (.A(_06725_),
    .X(_01092_));
 sky130_fd_sc_hd__mux2_1 _13322_ (.A0(_04992_),
    .A1(\regs[25][5] ),
    .S(_06720_),
    .X(_06726_));
 sky130_fd_sc_hd__clkbuf_1 _13323_ (.A(_06726_),
    .X(_01093_));
 sky130_fd_sc_hd__mux2_1 _13324_ (.A0(_05030_),
    .A1(\regs[25][6] ),
    .S(_06720_),
    .X(_06727_));
 sky130_fd_sc_hd__clkbuf_1 _13325_ (.A(_06727_),
    .X(_01094_));
 sky130_fd_sc_hd__mux2_1 _13326_ (.A0(_05080_),
    .A1(\regs[25][7] ),
    .S(_06720_),
    .X(_06728_));
 sky130_fd_sc_hd__clkbuf_1 _13327_ (.A(_06728_),
    .X(_01095_));
 sky130_fd_sc_hd__mux2_1 _13328_ (.A0(_05121_),
    .A1(\regs[25][8] ),
    .S(_06720_),
    .X(_06729_));
 sky130_fd_sc_hd__clkbuf_1 _13329_ (.A(_06729_),
    .X(_01096_));
 sky130_fd_sc_hd__mux2_1 _13330_ (.A0(_05157_),
    .A1(\regs[25][9] ),
    .S(_06720_),
    .X(_06730_));
 sky130_fd_sc_hd__clkbuf_1 _13331_ (.A(_06730_),
    .X(_01097_));
 sky130_fd_sc_hd__buf_6 _13332_ (.A(_06719_),
    .X(_06731_));
 sky130_fd_sc_hd__mux2_1 _13333_ (.A0(_05187_),
    .A1(\regs[25][10] ),
    .S(_06731_),
    .X(_06732_));
 sky130_fd_sc_hd__clkbuf_1 _13334_ (.A(_06732_),
    .X(_01098_));
 sky130_fd_sc_hd__mux2_1 _13335_ (.A0(_05224_),
    .A1(\regs[25][11] ),
    .S(_06731_),
    .X(_06733_));
 sky130_fd_sc_hd__clkbuf_1 _13336_ (.A(_06733_),
    .X(_01099_));
 sky130_fd_sc_hd__mux2_1 _13337_ (.A0(_05263_),
    .A1(\regs[25][12] ),
    .S(_06731_),
    .X(_06734_));
 sky130_fd_sc_hd__clkbuf_1 _13338_ (.A(_06734_),
    .X(_01100_));
 sky130_fd_sc_hd__mux2_1 _13339_ (.A0(_05296_),
    .A1(\regs[25][13] ),
    .S(_06731_),
    .X(_06735_));
 sky130_fd_sc_hd__clkbuf_1 _13340_ (.A(_06735_),
    .X(_01101_));
 sky130_fd_sc_hd__mux2_1 _13341_ (.A0(_05329_),
    .A1(\regs[25][14] ),
    .S(_06731_),
    .X(_06736_));
 sky130_fd_sc_hd__clkbuf_1 _13342_ (.A(_06736_),
    .X(_01102_));
 sky130_fd_sc_hd__mux2_1 _13343_ (.A0(_05359_),
    .A1(\regs[25][15] ),
    .S(_06731_),
    .X(_06737_));
 sky130_fd_sc_hd__clkbuf_1 _13344_ (.A(_06737_),
    .X(_01103_));
 sky130_fd_sc_hd__mux2_1 _13345_ (.A0(_05400_),
    .A1(\regs[25][16] ),
    .S(_06731_),
    .X(_06738_));
 sky130_fd_sc_hd__clkbuf_1 _13346_ (.A(_06738_),
    .X(_01104_));
 sky130_fd_sc_hd__mux2_1 _13347_ (.A0(_05424_),
    .A1(\regs[25][17] ),
    .S(_06731_),
    .X(_06739_));
 sky130_fd_sc_hd__clkbuf_1 _13348_ (.A(_06739_),
    .X(_01105_));
 sky130_fd_sc_hd__mux2_1 _13349_ (.A0(_05452_),
    .A1(\regs[25][18] ),
    .S(_06731_),
    .X(_06740_));
 sky130_fd_sc_hd__clkbuf_1 _13350_ (.A(_06740_),
    .X(_01106_));
 sky130_fd_sc_hd__mux2_1 _13351_ (.A0(_05477_),
    .A1(\regs[25][19] ),
    .S(_06731_),
    .X(_06741_));
 sky130_fd_sc_hd__clkbuf_1 _13352_ (.A(_06741_),
    .X(_01107_));
 sky130_fd_sc_hd__buf_4 _13353_ (.A(_06719_),
    .X(_06742_));
 sky130_fd_sc_hd__mux2_1 _13354_ (.A0(_05514_),
    .A1(\regs[25][20] ),
    .S(_06742_),
    .X(_06743_));
 sky130_fd_sc_hd__clkbuf_1 _13355_ (.A(_06743_),
    .X(_01108_));
 sky130_fd_sc_hd__mux2_1 _13356_ (.A0(_05541_),
    .A1(\regs[25][21] ),
    .S(_06742_),
    .X(_06744_));
 sky130_fd_sc_hd__clkbuf_1 _13357_ (.A(_06744_),
    .X(_01109_));
 sky130_fd_sc_hd__mux2_1 _13358_ (.A0(_05570_),
    .A1(\regs[25][22] ),
    .S(_06742_),
    .X(_06745_));
 sky130_fd_sc_hd__clkbuf_1 _13359_ (.A(_06745_),
    .X(_01110_));
 sky130_fd_sc_hd__mux2_1 _13360_ (.A0(_05600_),
    .A1(\regs[25][23] ),
    .S(_06742_),
    .X(_06746_));
 sky130_fd_sc_hd__clkbuf_1 _13361_ (.A(_06746_),
    .X(_01111_));
 sky130_fd_sc_hd__mux2_1 _13362_ (.A0(_05636_),
    .A1(\regs[25][24] ),
    .S(_06742_),
    .X(_06747_));
 sky130_fd_sc_hd__clkbuf_1 _13363_ (.A(_06747_),
    .X(_01112_));
 sky130_fd_sc_hd__mux2_1 _13364_ (.A0(_05660_),
    .A1(\regs[25][25] ),
    .S(_06742_),
    .X(_06748_));
 sky130_fd_sc_hd__clkbuf_1 _13365_ (.A(_06748_),
    .X(_01113_));
 sky130_fd_sc_hd__mux2_1 _13366_ (.A0(_05684_),
    .A1(\regs[25][26] ),
    .S(_06742_),
    .X(_06749_));
 sky130_fd_sc_hd__clkbuf_1 _13367_ (.A(_06749_),
    .X(_01114_));
 sky130_fd_sc_hd__mux2_1 _13368_ (.A0(_05708_),
    .A1(\regs[25][27] ),
    .S(_06742_),
    .X(_06750_));
 sky130_fd_sc_hd__clkbuf_1 _13369_ (.A(_06750_),
    .X(_01115_));
 sky130_fd_sc_hd__mux2_1 _13370_ (.A0(_05735_),
    .A1(\regs[25][28] ),
    .S(_06742_),
    .X(_06751_));
 sky130_fd_sc_hd__clkbuf_1 _13371_ (.A(_06751_),
    .X(_01116_));
 sky130_fd_sc_hd__mux2_1 _13372_ (.A0(_05763_),
    .A1(\regs[25][29] ),
    .S(_06742_),
    .X(_06752_));
 sky130_fd_sc_hd__clkbuf_1 _13373_ (.A(_06752_),
    .X(_01117_));
 sky130_fd_sc_hd__mux2_1 _13374_ (.A0(_05787_),
    .A1(\regs[25][30] ),
    .S(_06719_),
    .X(_06753_));
 sky130_fd_sc_hd__clkbuf_1 _13375_ (.A(_06753_),
    .X(_01118_));
 sky130_fd_sc_hd__mux2_1 _13376_ (.A0(_05811_),
    .A1(\regs[25][31] ),
    .S(_06719_),
    .X(_06754_));
 sky130_fd_sc_hd__clkbuf_1 _13377_ (.A(_06754_),
    .X(_01119_));
 sky130_fd_sc_hd__nand2_2 _13378_ (.A(_05884_),
    .B(_06682_),
    .Y(_06755_));
 sky130_fd_sc_hd__buf_4 _13379_ (.A(_06755_),
    .X(_06756_));
 sky130_fd_sc_hd__mux2_1 _13380_ (.A0(_04762_),
    .A1(\regs[26][0] ),
    .S(_06756_),
    .X(_06757_));
 sky130_fd_sc_hd__clkbuf_1 _13381_ (.A(_06757_),
    .X(_01120_));
 sky130_fd_sc_hd__mux2_1 _13382_ (.A0(_04818_),
    .A1(\regs[26][1] ),
    .S(_06756_),
    .X(_06758_));
 sky130_fd_sc_hd__clkbuf_1 _13383_ (.A(_06758_),
    .X(_01121_));
 sky130_fd_sc_hd__mux2_1 _13384_ (.A0(_04858_),
    .A1(\regs[26][2] ),
    .S(_06756_),
    .X(_06759_));
 sky130_fd_sc_hd__clkbuf_1 _13385_ (.A(_06759_),
    .X(_01122_));
 sky130_fd_sc_hd__mux2_1 _13386_ (.A0(_04904_),
    .A1(\regs[26][3] ),
    .S(_06756_),
    .X(_06760_));
 sky130_fd_sc_hd__clkbuf_1 _13387_ (.A(_06760_),
    .X(_01123_));
 sky130_fd_sc_hd__mux2_1 _13388_ (.A0(_04952_),
    .A1(\regs[26][4] ),
    .S(_06756_),
    .X(_06761_));
 sky130_fd_sc_hd__clkbuf_1 _13389_ (.A(_06761_),
    .X(_01124_));
 sky130_fd_sc_hd__mux2_1 _13390_ (.A0(_04992_),
    .A1(\regs[26][5] ),
    .S(_06756_),
    .X(_06762_));
 sky130_fd_sc_hd__clkbuf_1 _13391_ (.A(_06762_),
    .X(_01125_));
 sky130_fd_sc_hd__mux2_1 _13392_ (.A0(_05030_),
    .A1(\regs[26][6] ),
    .S(_06756_),
    .X(_06763_));
 sky130_fd_sc_hd__clkbuf_1 _13393_ (.A(_06763_),
    .X(_01126_));
 sky130_fd_sc_hd__mux2_1 _13394_ (.A0(_05080_),
    .A1(\regs[26][7] ),
    .S(_06756_),
    .X(_06764_));
 sky130_fd_sc_hd__clkbuf_1 _13395_ (.A(_06764_),
    .X(_01127_));
 sky130_fd_sc_hd__mux2_1 _13396_ (.A0(_05121_),
    .A1(\regs[26][8] ),
    .S(_06756_),
    .X(_06765_));
 sky130_fd_sc_hd__clkbuf_1 _13397_ (.A(_06765_),
    .X(_01128_));
 sky130_fd_sc_hd__mux2_1 _13398_ (.A0(_05157_),
    .A1(\regs[26][9] ),
    .S(_06756_),
    .X(_06766_));
 sky130_fd_sc_hd__clkbuf_1 _13399_ (.A(_06766_),
    .X(_01129_));
 sky130_fd_sc_hd__clkbuf_8 _13400_ (.A(_06755_),
    .X(_06767_));
 sky130_fd_sc_hd__mux2_1 _13401_ (.A0(_05187_),
    .A1(\regs[26][10] ),
    .S(_06767_),
    .X(_06768_));
 sky130_fd_sc_hd__clkbuf_1 _13402_ (.A(_06768_),
    .X(_01130_));
 sky130_fd_sc_hd__mux2_1 _13403_ (.A0(_05224_),
    .A1(\regs[26][11] ),
    .S(_06767_),
    .X(_06769_));
 sky130_fd_sc_hd__clkbuf_1 _13404_ (.A(_06769_),
    .X(_01131_));
 sky130_fd_sc_hd__mux2_1 _13405_ (.A0(_05263_),
    .A1(\regs[26][12] ),
    .S(_06767_),
    .X(_06770_));
 sky130_fd_sc_hd__clkbuf_1 _13406_ (.A(_06770_),
    .X(_01132_));
 sky130_fd_sc_hd__mux2_1 _13407_ (.A0(_05296_),
    .A1(\regs[26][13] ),
    .S(_06767_),
    .X(_06771_));
 sky130_fd_sc_hd__clkbuf_1 _13408_ (.A(_06771_),
    .X(_01133_));
 sky130_fd_sc_hd__mux2_1 _13409_ (.A0(_05329_),
    .A1(\regs[26][14] ),
    .S(_06767_),
    .X(_06772_));
 sky130_fd_sc_hd__clkbuf_1 _13410_ (.A(_06772_),
    .X(_01134_));
 sky130_fd_sc_hd__mux2_1 _13411_ (.A0(_05359_),
    .A1(\regs[26][15] ),
    .S(_06767_),
    .X(_06773_));
 sky130_fd_sc_hd__clkbuf_1 _13412_ (.A(_06773_),
    .X(_01135_));
 sky130_fd_sc_hd__mux2_1 _13413_ (.A0(_05400_),
    .A1(\regs[26][16] ),
    .S(_06767_),
    .X(_06774_));
 sky130_fd_sc_hd__clkbuf_1 _13414_ (.A(_06774_),
    .X(_01136_));
 sky130_fd_sc_hd__mux2_1 _13415_ (.A0(_05424_),
    .A1(\regs[26][17] ),
    .S(_06767_),
    .X(_06775_));
 sky130_fd_sc_hd__clkbuf_1 _13416_ (.A(_06775_),
    .X(_01137_));
 sky130_fd_sc_hd__mux2_1 _13417_ (.A0(_05452_),
    .A1(\regs[26][18] ),
    .S(_06767_),
    .X(_06776_));
 sky130_fd_sc_hd__clkbuf_1 _13418_ (.A(_06776_),
    .X(_01138_));
 sky130_fd_sc_hd__mux2_1 _13419_ (.A0(_05477_),
    .A1(\regs[26][19] ),
    .S(_06767_),
    .X(_06777_));
 sky130_fd_sc_hd__clkbuf_1 _13420_ (.A(_06777_),
    .X(_01139_));
 sky130_fd_sc_hd__buf_4 _13421_ (.A(_06755_),
    .X(_06778_));
 sky130_fd_sc_hd__mux2_1 _13422_ (.A0(_05514_),
    .A1(\regs[26][20] ),
    .S(_06778_),
    .X(_06779_));
 sky130_fd_sc_hd__clkbuf_1 _13423_ (.A(_06779_),
    .X(_01140_));
 sky130_fd_sc_hd__mux2_1 _13424_ (.A0(_05541_),
    .A1(\regs[26][21] ),
    .S(_06778_),
    .X(_06780_));
 sky130_fd_sc_hd__clkbuf_1 _13425_ (.A(_06780_),
    .X(_01141_));
 sky130_fd_sc_hd__mux2_1 _13426_ (.A0(_05570_),
    .A1(\regs[26][22] ),
    .S(_06778_),
    .X(_06781_));
 sky130_fd_sc_hd__clkbuf_1 _13427_ (.A(_06781_),
    .X(_01142_));
 sky130_fd_sc_hd__mux2_1 _13428_ (.A0(_05600_),
    .A1(\regs[26][23] ),
    .S(_06778_),
    .X(_06782_));
 sky130_fd_sc_hd__clkbuf_1 _13429_ (.A(_06782_),
    .X(_01143_));
 sky130_fd_sc_hd__mux2_1 _13430_ (.A0(_05636_),
    .A1(\regs[26][24] ),
    .S(_06778_),
    .X(_06783_));
 sky130_fd_sc_hd__clkbuf_1 _13431_ (.A(_06783_),
    .X(_01144_));
 sky130_fd_sc_hd__mux2_1 _13432_ (.A0(_05660_),
    .A1(\regs[26][25] ),
    .S(_06778_),
    .X(_06784_));
 sky130_fd_sc_hd__clkbuf_1 _13433_ (.A(_06784_),
    .X(_01145_));
 sky130_fd_sc_hd__mux2_1 _13434_ (.A0(_05684_),
    .A1(\regs[26][26] ),
    .S(_06778_),
    .X(_06785_));
 sky130_fd_sc_hd__clkbuf_1 _13435_ (.A(_06785_),
    .X(_01146_));
 sky130_fd_sc_hd__mux2_1 _13436_ (.A0(_05708_),
    .A1(\regs[26][27] ),
    .S(_06778_),
    .X(_06786_));
 sky130_fd_sc_hd__clkbuf_1 _13437_ (.A(_06786_),
    .X(_01147_));
 sky130_fd_sc_hd__mux2_1 _13438_ (.A0(_05735_),
    .A1(\regs[26][28] ),
    .S(_06778_),
    .X(_06787_));
 sky130_fd_sc_hd__clkbuf_1 _13439_ (.A(_06787_),
    .X(_01148_));
 sky130_fd_sc_hd__mux2_1 _13440_ (.A0(_05763_),
    .A1(\regs[26][29] ),
    .S(_06778_),
    .X(_06788_));
 sky130_fd_sc_hd__clkbuf_1 _13441_ (.A(_06788_),
    .X(_01149_));
 sky130_fd_sc_hd__mux2_1 _13442_ (.A0(_05787_),
    .A1(\regs[26][30] ),
    .S(_06755_),
    .X(_06789_));
 sky130_fd_sc_hd__clkbuf_1 _13443_ (.A(_06789_),
    .X(_01150_));
 sky130_fd_sc_hd__mux2_1 _13444_ (.A0(_05811_),
    .A1(\regs[26][31] ),
    .S(_06755_),
    .X(_06790_));
 sky130_fd_sc_hd__clkbuf_1 _13445_ (.A(_06790_),
    .X(_01151_));
 sky130_fd_sc_hd__and2_2 _13446_ (.A(_05815_),
    .B(_05884_),
    .X(_06791_));
 sky130_fd_sc_hd__buf_6 _13447_ (.A(_06791_),
    .X(_06792_));
 sky130_fd_sc_hd__mux2_1 _13448_ (.A0(\regs[6][0] ),
    .A1(_06291_),
    .S(_06792_),
    .X(_06793_));
 sky130_fd_sc_hd__clkbuf_1 _13449_ (.A(_06793_),
    .X(_01152_));
 sky130_fd_sc_hd__mux2_1 _13450_ (.A0(\regs[6][1] ),
    .A1(_06295_),
    .S(_06792_),
    .X(_06794_));
 sky130_fd_sc_hd__clkbuf_1 _13451_ (.A(_06794_),
    .X(_01153_));
 sky130_fd_sc_hd__mux2_1 _13452_ (.A0(\regs[6][2] ),
    .A1(_06297_),
    .S(_06792_),
    .X(_06795_));
 sky130_fd_sc_hd__clkbuf_1 _13453_ (.A(_06795_),
    .X(_01154_));
 sky130_fd_sc_hd__mux2_1 _13454_ (.A0(\regs[6][3] ),
    .A1(_06299_),
    .S(_06792_),
    .X(_06796_));
 sky130_fd_sc_hd__clkbuf_1 _13455_ (.A(_06796_),
    .X(_01155_));
 sky130_fd_sc_hd__mux2_1 _13456_ (.A0(\regs[6][4] ),
    .A1(_06301_),
    .S(_06792_),
    .X(_06797_));
 sky130_fd_sc_hd__clkbuf_1 _13457_ (.A(_06797_),
    .X(_01156_));
 sky130_fd_sc_hd__mux2_1 _13458_ (.A0(\regs[6][5] ),
    .A1(_06303_),
    .S(_06792_),
    .X(_06798_));
 sky130_fd_sc_hd__clkbuf_1 _13459_ (.A(_06798_),
    .X(_01157_));
 sky130_fd_sc_hd__mux2_1 _13460_ (.A0(\regs[6][6] ),
    .A1(_06305_),
    .S(_06792_),
    .X(_06799_));
 sky130_fd_sc_hd__clkbuf_1 _13461_ (.A(_06799_),
    .X(_01158_));
 sky130_fd_sc_hd__mux2_1 _13462_ (.A0(\regs[6][7] ),
    .A1(_06307_),
    .S(_06792_),
    .X(_06800_));
 sky130_fd_sc_hd__clkbuf_1 _13463_ (.A(_06800_),
    .X(_01159_));
 sky130_fd_sc_hd__mux2_1 _13464_ (.A0(\regs[6][8] ),
    .A1(_06309_),
    .S(_06792_),
    .X(_06801_));
 sky130_fd_sc_hd__clkbuf_1 _13465_ (.A(_06801_),
    .X(_01160_));
 sky130_fd_sc_hd__mux2_1 _13466_ (.A0(\regs[6][9] ),
    .A1(_06311_),
    .S(_06792_),
    .X(_06802_));
 sky130_fd_sc_hd__clkbuf_1 _13467_ (.A(_06802_),
    .X(_01161_));
 sky130_fd_sc_hd__buf_4 _13468_ (.A(_06791_),
    .X(_06803_));
 sky130_fd_sc_hd__mux2_1 _13469_ (.A0(\regs[6][10] ),
    .A1(_06313_),
    .S(_06803_),
    .X(_06804_));
 sky130_fd_sc_hd__clkbuf_1 _13470_ (.A(_06804_),
    .X(_01162_));
 sky130_fd_sc_hd__mux2_1 _13471_ (.A0(\regs[6][11] ),
    .A1(_06316_),
    .S(_06803_),
    .X(_06805_));
 sky130_fd_sc_hd__clkbuf_1 _13472_ (.A(_06805_),
    .X(_01163_));
 sky130_fd_sc_hd__mux2_1 _13473_ (.A0(\regs[6][12] ),
    .A1(_06318_),
    .S(_06803_),
    .X(_06806_));
 sky130_fd_sc_hd__clkbuf_1 _13474_ (.A(_06806_),
    .X(_01164_));
 sky130_fd_sc_hd__mux2_1 _13475_ (.A0(\regs[6][13] ),
    .A1(_06320_),
    .S(_06803_),
    .X(_06807_));
 sky130_fd_sc_hd__clkbuf_1 _13476_ (.A(_06807_),
    .X(_01165_));
 sky130_fd_sc_hd__mux2_1 _13477_ (.A0(\regs[6][14] ),
    .A1(_06322_),
    .S(_06803_),
    .X(_06808_));
 sky130_fd_sc_hd__clkbuf_1 _13478_ (.A(_06808_),
    .X(_01166_));
 sky130_fd_sc_hd__mux2_1 _13479_ (.A0(\regs[6][15] ),
    .A1(_06324_),
    .S(_06803_),
    .X(_06809_));
 sky130_fd_sc_hd__clkbuf_1 _13480_ (.A(_06809_),
    .X(_01167_));
 sky130_fd_sc_hd__mux2_1 _13481_ (.A0(\regs[6][16] ),
    .A1(_06326_),
    .S(_06803_),
    .X(_06810_));
 sky130_fd_sc_hd__clkbuf_1 _13482_ (.A(_06810_),
    .X(_01168_));
 sky130_fd_sc_hd__mux2_1 _13483_ (.A0(\regs[6][17] ),
    .A1(_06328_),
    .S(_06803_),
    .X(_06811_));
 sky130_fd_sc_hd__clkbuf_1 _13484_ (.A(_06811_),
    .X(_01169_));
 sky130_fd_sc_hd__mux2_1 _13485_ (.A0(\regs[6][18] ),
    .A1(_06330_),
    .S(_06803_),
    .X(_06812_));
 sky130_fd_sc_hd__clkbuf_1 _13486_ (.A(_06812_),
    .X(_01170_));
 sky130_fd_sc_hd__mux2_1 _13487_ (.A0(\regs[6][19] ),
    .A1(_06332_),
    .S(_06803_),
    .X(_06813_));
 sky130_fd_sc_hd__clkbuf_1 _13488_ (.A(_06813_),
    .X(_01171_));
 sky130_fd_sc_hd__buf_6 _13489_ (.A(_06791_),
    .X(_06814_));
 sky130_fd_sc_hd__mux2_1 _13490_ (.A0(\regs[6][20] ),
    .A1(_06334_),
    .S(_06814_),
    .X(_06815_));
 sky130_fd_sc_hd__clkbuf_1 _13491_ (.A(_06815_),
    .X(_01172_));
 sky130_fd_sc_hd__mux2_1 _13492_ (.A0(\regs[6][21] ),
    .A1(_06337_),
    .S(_06814_),
    .X(_06816_));
 sky130_fd_sc_hd__clkbuf_1 _13493_ (.A(_06816_),
    .X(_01173_));
 sky130_fd_sc_hd__mux2_1 _13494_ (.A0(\regs[6][22] ),
    .A1(_06339_),
    .S(_06814_),
    .X(_06817_));
 sky130_fd_sc_hd__clkbuf_1 _13495_ (.A(_06817_),
    .X(_01174_));
 sky130_fd_sc_hd__mux2_1 _13496_ (.A0(\regs[6][23] ),
    .A1(_06341_),
    .S(_06814_),
    .X(_06818_));
 sky130_fd_sc_hd__clkbuf_1 _13497_ (.A(_06818_),
    .X(_01175_));
 sky130_fd_sc_hd__mux2_1 _13498_ (.A0(\regs[6][24] ),
    .A1(_06343_),
    .S(_06814_),
    .X(_06819_));
 sky130_fd_sc_hd__clkbuf_1 _13499_ (.A(_06819_),
    .X(_01176_));
 sky130_fd_sc_hd__mux2_1 _13500_ (.A0(\regs[6][25] ),
    .A1(_06345_),
    .S(_06814_),
    .X(_06820_));
 sky130_fd_sc_hd__clkbuf_1 _13501_ (.A(_06820_),
    .X(_01177_));
 sky130_fd_sc_hd__mux2_1 _13502_ (.A0(\regs[6][26] ),
    .A1(_06347_),
    .S(_06814_),
    .X(_06821_));
 sky130_fd_sc_hd__clkbuf_1 _13503_ (.A(_06821_),
    .X(_01178_));
 sky130_fd_sc_hd__mux2_1 _13504_ (.A0(\regs[6][27] ),
    .A1(_06349_),
    .S(_06814_),
    .X(_06822_));
 sky130_fd_sc_hd__clkbuf_1 _13505_ (.A(_06822_),
    .X(_01179_));
 sky130_fd_sc_hd__mux2_1 _13506_ (.A0(\regs[6][28] ),
    .A1(_06351_),
    .S(_06814_),
    .X(_06823_));
 sky130_fd_sc_hd__clkbuf_1 _13507_ (.A(_06823_),
    .X(_01180_));
 sky130_fd_sc_hd__mux2_1 _13508_ (.A0(\regs[6][29] ),
    .A1(_06353_),
    .S(_06814_),
    .X(_06824_));
 sky130_fd_sc_hd__clkbuf_1 _13509_ (.A(_06824_),
    .X(_01181_));
 sky130_fd_sc_hd__mux2_1 _13510_ (.A0(\regs[6][30] ),
    .A1(_06355_),
    .S(_06791_),
    .X(_06825_));
 sky130_fd_sc_hd__clkbuf_1 _13511_ (.A(_06825_),
    .X(_01182_));
 sky130_fd_sc_hd__mux2_1 _13512_ (.A0(\regs[6][31] ),
    .A1(_06357_),
    .S(_06791_),
    .X(_06826_));
 sky130_fd_sc_hd__clkbuf_1 _13513_ (.A(_06826_),
    .X(_01183_));
 sky130_fd_sc_hd__nand2_2 _13514_ (.A(_05814_),
    .B(_06682_),
    .Y(_06827_));
 sky130_fd_sc_hd__buf_4 _13515_ (.A(_06827_),
    .X(_06828_));
 sky130_fd_sc_hd__mux2_1 _13516_ (.A0(_04762_),
    .A1(\regs[27][0] ),
    .S(_06828_),
    .X(_06829_));
 sky130_fd_sc_hd__clkbuf_1 _13517_ (.A(_06829_),
    .X(_01184_));
 sky130_fd_sc_hd__mux2_1 _13518_ (.A0(_04818_),
    .A1(\regs[27][1] ),
    .S(_06828_),
    .X(_06830_));
 sky130_fd_sc_hd__clkbuf_1 _13519_ (.A(_06830_),
    .X(_01185_));
 sky130_fd_sc_hd__mux2_1 _13520_ (.A0(_04858_),
    .A1(\regs[27][2] ),
    .S(_06828_),
    .X(_06831_));
 sky130_fd_sc_hd__clkbuf_1 _13521_ (.A(_06831_),
    .X(_01186_));
 sky130_fd_sc_hd__mux2_1 _13522_ (.A0(_04904_),
    .A1(\regs[27][3] ),
    .S(_06828_),
    .X(_06832_));
 sky130_fd_sc_hd__clkbuf_1 _13523_ (.A(_06832_),
    .X(_01187_));
 sky130_fd_sc_hd__mux2_1 _13524_ (.A0(_04952_),
    .A1(\regs[27][4] ),
    .S(_06828_),
    .X(_06833_));
 sky130_fd_sc_hd__clkbuf_1 _13525_ (.A(_06833_),
    .X(_01188_));
 sky130_fd_sc_hd__mux2_1 _13526_ (.A0(_04992_),
    .A1(\regs[27][5] ),
    .S(_06828_),
    .X(_06834_));
 sky130_fd_sc_hd__clkbuf_1 _13527_ (.A(_06834_),
    .X(_01189_));
 sky130_fd_sc_hd__mux2_1 _13528_ (.A0(_05030_),
    .A1(\regs[27][6] ),
    .S(_06828_),
    .X(_06835_));
 sky130_fd_sc_hd__clkbuf_1 _13529_ (.A(_06835_),
    .X(_01190_));
 sky130_fd_sc_hd__mux2_1 _13530_ (.A0(_05080_),
    .A1(\regs[27][7] ),
    .S(_06828_),
    .X(_06836_));
 sky130_fd_sc_hd__clkbuf_1 _13531_ (.A(_06836_),
    .X(_01191_));
 sky130_fd_sc_hd__mux2_1 _13532_ (.A0(_05121_),
    .A1(\regs[27][8] ),
    .S(_06828_),
    .X(_06837_));
 sky130_fd_sc_hd__clkbuf_1 _13533_ (.A(_06837_),
    .X(_01192_));
 sky130_fd_sc_hd__mux2_1 _13534_ (.A0(_05157_),
    .A1(\regs[27][9] ),
    .S(_06828_),
    .X(_06838_));
 sky130_fd_sc_hd__clkbuf_1 _13535_ (.A(_06838_),
    .X(_01193_));
 sky130_fd_sc_hd__clkbuf_8 _13536_ (.A(_06827_),
    .X(_06839_));
 sky130_fd_sc_hd__mux2_1 _13537_ (.A0(_05187_),
    .A1(\regs[27][10] ),
    .S(_06839_),
    .X(_06840_));
 sky130_fd_sc_hd__clkbuf_1 _13538_ (.A(_06840_),
    .X(_01194_));
 sky130_fd_sc_hd__mux2_1 _13539_ (.A0(_05224_),
    .A1(\regs[27][11] ),
    .S(_06839_),
    .X(_06841_));
 sky130_fd_sc_hd__clkbuf_1 _13540_ (.A(_06841_),
    .X(_01195_));
 sky130_fd_sc_hd__mux2_1 _13541_ (.A0(_05263_),
    .A1(\regs[27][12] ),
    .S(_06839_),
    .X(_06842_));
 sky130_fd_sc_hd__clkbuf_1 _13542_ (.A(_06842_),
    .X(_01196_));
 sky130_fd_sc_hd__mux2_1 _13543_ (.A0(_05296_),
    .A1(\regs[27][13] ),
    .S(_06839_),
    .X(_06843_));
 sky130_fd_sc_hd__clkbuf_1 _13544_ (.A(_06843_),
    .X(_01197_));
 sky130_fd_sc_hd__mux2_1 _13545_ (.A0(_05329_),
    .A1(\regs[27][14] ),
    .S(_06839_),
    .X(_06844_));
 sky130_fd_sc_hd__clkbuf_1 _13546_ (.A(_06844_),
    .X(_01198_));
 sky130_fd_sc_hd__mux2_1 _13547_ (.A0(_05359_),
    .A1(\regs[27][15] ),
    .S(_06839_),
    .X(_06845_));
 sky130_fd_sc_hd__clkbuf_1 _13548_ (.A(_06845_),
    .X(_01199_));
 sky130_fd_sc_hd__mux2_1 _13549_ (.A0(_05400_),
    .A1(\regs[27][16] ),
    .S(_06839_),
    .X(_06846_));
 sky130_fd_sc_hd__clkbuf_1 _13550_ (.A(_06846_),
    .X(_01200_));
 sky130_fd_sc_hd__mux2_1 _13551_ (.A0(_05424_),
    .A1(\regs[27][17] ),
    .S(_06839_),
    .X(_06847_));
 sky130_fd_sc_hd__clkbuf_1 _13552_ (.A(_06847_),
    .X(_01201_));
 sky130_fd_sc_hd__mux2_1 _13553_ (.A0(_05452_),
    .A1(\regs[27][18] ),
    .S(_06839_),
    .X(_06848_));
 sky130_fd_sc_hd__clkbuf_1 _13554_ (.A(_06848_),
    .X(_01202_));
 sky130_fd_sc_hd__mux2_1 _13555_ (.A0(_05477_),
    .A1(\regs[27][19] ),
    .S(_06839_),
    .X(_06849_));
 sky130_fd_sc_hd__clkbuf_1 _13556_ (.A(_06849_),
    .X(_01203_));
 sky130_fd_sc_hd__buf_4 _13557_ (.A(_06827_),
    .X(_06850_));
 sky130_fd_sc_hd__mux2_1 _13558_ (.A0(_05514_),
    .A1(\regs[27][20] ),
    .S(_06850_),
    .X(_06851_));
 sky130_fd_sc_hd__clkbuf_1 _13559_ (.A(_06851_),
    .X(_01204_));
 sky130_fd_sc_hd__mux2_1 _13560_ (.A0(_05541_),
    .A1(\regs[27][21] ),
    .S(_06850_),
    .X(_06852_));
 sky130_fd_sc_hd__clkbuf_1 _13561_ (.A(_06852_),
    .X(_01205_));
 sky130_fd_sc_hd__mux2_1 _13562_ (.A0(_05570_),
    .A1(\regs[27][22] ),
    .S(_06850_),
    .X(_06853_));
 sky130_fd_sc_hd__clkbuf_1 _13563_ (.A(_06853_),
    .X(_01206_));
 sky130_fd_sc_hd__mux2_1 _13564_ (.A0(_05600_),
    .A1(\regs[27][23] ),
    .S(_06850_),
    .X(_06854_));
 sky130_fd_sc_hd__clkbuf_1 _13565_ (.A(_06854_),
    .X(_01207_));
 sky130_fd_sc_hd__mux2_1 _13566_ (.A0(_05636_),
    .A1(\regs[27][24] ),
    .S(_06850_),
    .X(_06855_));
 sky130_fd_sc_hd__clkbuf_1 _13567_ (.A(_06855_),
    .X(_01208_));
 sky130_fd_sc_hd__mux2_1 _13568_ (.A0(_05660_),
    .A1(\regs[27][25] ),
    .S(_06850_),
    .X(_06856_));
 sky130_fd_sc_hd__clkbuf_1 _13569_ (.A(_06856_),
    .X(_01209_));
 sky130_fd_sc_hd__mux2_1 _13570_ (.A0(_05684_),
    .A1(\regs[27][26] ),
    .S(_06850_),
    .X(_06857_));
 sky130_fd_sc_hd__clkbuf_1 _13571_ (.A(_06857_),
    .X(_01210_));
 sky130_fd_sc_hd__mux2_1 _13572_ (.A0(_05708_),
    .A1(\regs[27][27] ),
    .S(_06850_),
    .X(_06858_));
 sky130_fd_sc_hd__clkbuf_1 _13573_ (.A(_06858_),
    .X(_01211_));
 sky130_fd_sc_hd__mux2_1 _13574_ (.A0(_05735_),
    .A1(\regs[27][28] ),
    .S(_06850_),
    .X(_06859_));
 sky130_fd_sc_hd__clkbuf_1 _13575_ (.A(_06859_),
    .X(_01212_));
 sky130_fd_sc_hd__mux2_1 _13576_ (.A0(_05763_),
    .A1(\regs[27][29] ),
    .S(_06850_),
    .X(_06860_));
 sky130_fd_sc_hd__clkbuf_1 _13577_ (.A(_06860_),
    .X(_01213_));
 sky130_fd_sc_hd__mux2_1 _13578_ (.A0(_05787_),
    .A1(\regs[27][30] ),
    .S(_06827_),
    .X(_06861_));
 sky130_fd_sc_hd__clkbuf_1 _13579_ (.A(_06861_),
    .X(_01214_));
 sky130_fd_sc_hd__mux2_1 _13580_ (.A0(_05811_),
    .A1(\regs[27][31] ),
    .S(_06827_),
    .X(_06862_));
 sky130_fd_sc_hd__clkbuf_1 _13581_ (.A(_06862_),
    .X(_01215_));
 sky130_fd_sc_hd__nor2_2 _13582_ (.A(_04758_),
    .B(_06218_),
    .Y(_06863_));
 sky130_fd_sc_hd__buf_6 _13583_ (.A(_06863_),
    .X(_06864_));
 sky130_fd_sc_hd__mux2_1 _13584_ (.A0(\regs[28][0] ),
    .A1(_06291_),
    .S(_06864_),
    .X(_06865_));
 sky130_fd_sc_hd__clkbuf_1 _13585_ (.A(_06865_),
    .X(_01216_));
 sky130_fd_sc_hd__mux2_1 _13586_ (.A0(\regs[28][1] ),
    .A1(_06295_),
    .S(_06864_),
    .X(_06866_));
 sky130_fd_sc_hd__clkbuf_1 _13587_ (.A(_06866_),
    .X(_01217_));
 sky130_fd_sc_hd__mux2_1 _13588_ (.A0(\regs[28][2] ),
    .A1(_06297_),
    .S(_06864_),
    .X(_06867_));
 sky130_fd_sc_hd__clkbuf_1 _13589_ (.A(_06867_),
    .X(_01218_));
 sky130_fd_sc_hd__mux2_1 _13590_ (.A0(\regs[28][3] ),
    .A1(_06299_),
    .S(_06864_),
    .X(_06868_));
 sky130_fd_sc_hd__clkbuf_1 _13591_ (.A(_06868_),
    .X(_01219_));
 sky130_fd_sc_hd__mux2_1 _13592_ (.A0(\regs[28][4] ),
    .A1(_06301_),
    .S(_06864_),
    .X(_06869_));
 sky130_fd_sc_hd__clkbuf_1 _13593_ (.A(_06869_),
    .X(_01220_));
 sky130_fd_sc_hd__mux2_1 _13594_ (.A0(\regs[28][5] ),
    .A1(_06303_),
    .S(_06864_),
    .X(_06870_));
 sky130_fd_sc_hd__clkbuf_1 _13595_ (.A(_06870_),
    .X(_01221_));
 sky130_fd_sc_hd__mux2_1 _13596_ (.A0(\regs[28][6] ),
    .A1(_06305_),
    .S(_06864_),
    .X(_06871_));
 sky130_fd_sc_hd__clkbuf_1 _13597_ (.A(_06871_),
    .X(_01222_));
 sky130_fd_sc_hd__mux2_1 _13598_ (.A0(\regs[28][7] ),
    .A1(_06307_),
    .S(_06864_),
    .X(_06872_));
 sky130_fd_sc_hd__clkbuf_1 _13599_ (.A(_06872_),
    .X(_01223_));
 sky130_fd_sc_hd__mux2_1 _13600_ (.A0(\regs[28][8] ),
    .A1(_06309_),
    .S(_06864_),
    .X(_06873_));
 sky130_fd_sc_hd__clkbuf_1 _13601_ (.A(_06873_),
    .X(_01224_));
 sky130_fd_sc_hd__mux2_1 _13602_ (.A0(\regs[28][9] ),
    .A1(_06311_),
    .S(_06864_),
    .X(_06874_));
 sky130_fd_sc_hd__clkbuf_1 _13603_ (.A(_06874_),
    .X(_01225_));
 sky130_fd_sc_hd__buf_4 _13604_ (.A(_06863_),
    .X(_06875_));
 sky130_fd_sc_hd__mux2_1 _13605_ (.A0(\regs[28][10] ),
    .A1(_06313_),
    .S(_06875_),
    .X(_06876_));
 sky130_fd_sc_hd__clkbuf_1 _13606_ (.A(_06876_),
    .X(_01226_));
 sky130_fd_sc_hd__mux2_1 _13607_ (.A0(\regs[28][11] ),
    .A1(_06316_),
    .S(_06875_),
    .X(_06877_));
 sky130_fd_sc_hd__clkbuf_1 _13608_ (.A(_06877_),
    .X(_01227_));
 sky130_fd_sc_hd__mux2_1 _13609_ (.A0(\regs[28][12] ),
    .A1(_06318_),
    .S(_06875_),
    .X(_06878_));
 sky130_fd_sc_hd__clkbuf_1 _13610_ (.A(_06878_),
    .X(_01228_));
 sky130_fd_sc_hd__mux2_1 _13611_ (.A0(\regs[28][13] ),
    .A1(_06320_),
    .S(_06875_),
    .X(_06879_));
 sky130_fd_sc_hd__clkbuf_1 _13612_ (.A(_06879_),
    .X(_01229_));
 sky130_fd_sc_hd__mux2_1 _13613_ (.A0(\regs[28][14] ),
    .A1(_06322_),
    .S(_06875_),
    .X(_06880_));
 sky130_fd_sc_hd__clkbuf_1 _13614_ (.A(_06880_),
    .X(_01230_));
 sky130_fd_sc_hd__mux2_1 _13615_ (.A0(\regs[28][15] ),
    .A1(_06324_),
    .S(_06875_),
    .X(_06881_));
 sky130_fd_sc_hd__clkbuf_1 _13616_ (.A(_06881_),
    .X(_01231_));
 sky130_fd_sc_hd__mux2_1 _13617_ (.A0(\regs[28][16] ),
    .A1(_06326_),
    .S(_06875_),
    .X(_06882_));
 sky130_fd_sc_hd__clkbuf_1 _13618_ (.A(_06882_),
    .X(_01232_));
 sky130_fd_sc_hd__mux2_1 _13619_ (.A0(\regs[28][17] ),
    .A1(_06328_),
    .S(_06875_),
    .X(_06883_));
 sky130_fd_sc_hd__clkbuf_1 _13620_ (.A(_06883_),
    .X(_01233_));
 sky130_fd_sc_hd__mux2_1 _13621_ (.A0(\regs[28][18] ),
    .A1(_06330_),
    .S(_06875_),
    .X(_06884_));
 sky130_fd_sc_hd__clkbuf_1 _13622_ (.A(_06884_),
    .X(_01234_));
 sky130_fd_sc_hd__mux2_1 _13623_ (.A0(\regs[28][19] ),
    .A1(_06332_),
    .S(_06875_),
    .X(_06885_));
 sky130_fd_sc_hd__clkbuf_1 _13624_ (.A(_06885_),
    .X(_01235_));
 sky130_fd_sc_hd__buf_4 _13625_ (.A(_06863_),
    .X(_06886_));
 sky130_fd_sc_hd__mux2_1 _13626_ (.A0(\regs[28][20] ),
    .A1(_06334_),
    .S(_06886_),
    .X(_06887_));
 sky130_fd_sc_hd__clkbuf_1 _13627_ (.A(_06887_),
    .X(_01236_));
 sky130_fd_sc_hd__mux2_1 _13628_ (.A0(\regs[28][21] ),
    .A1(_06337_),
    .S(_06886_),
    .X(_06888_));
 sky130_fd_sc_hd__clkbuf_1 _13629_ (.A(_06888_),
    .X(_01237_));
 sky130_fd_sc_hd__mux2_1 _13630_ (.A0(\regs[28][22] ),
    .A1(_06339_),
    .S(_06886_),
    .X(_06889_));
 sky130_fd_sc_hd__clkbuf_1 _13631_ (.A(_06889_),
    .X(_01238_));
 sky130_fd_sc_hd__mux2_1 _13632_ (.A0(\regs[28][23] ),
    .A1(_06341_),
    .S(_06886_),
    .X(_06890_));
 sky130_fd_sc_hd__clkbuf_1 _13633_ (.A(_06890_),
    .X(_01239_));
 sky130_fd_sc_hd__mux2_1 _13634_ (.A0(\regs[28][24] ),
    .A1(_06343_),
    .S(_06886_),
    .X(_06891_));
 sky130_fd_sc_hd__clkbuf_1 _13635_ (.A(_06891_),
    .X(_01240_));
 sky130_fd_sc_hd__mux2_1 _13636_ (.A0(\regs[28][25] ),
    .A1(_06345_),
    .S(_06886_),
    .X(_06892_));
 sky130_fd_sc_hd__clkbuf_1 _13637_ (.A(_06892_),
    .X(_01241_));
 sky130_fd_sc_hd__mux2_1 _13638_ (.A0(\regs[28][26] ),
    .A1(_06347_),
    .S(_06886_),
    .X(_06893_));
 sky130_fd_sc_hd__clkbuf_1 _13639_ (.A(_06893_),
    .X(_01242_));
 sky130_fd_sc_hd__mux2_1 _13640_ (.A0(\regs[28][27] ),
    .A1(_06349_),
    .S(_06886_),
    .X(_06894_));
 sky130_fd_sc_hd__clkbuf_1 _13641_ (.A(_06894_),
    .X(_01243_));
 sky130_fd_sc_hd__mux2_1 _13642_ (.A0(\regs[28][28] ),
    .A1(_06351_),
    .S(_06886_),
    .X(_06895_));
 sky130_fd_sc_hd__clkbuf_1 _13643_ (.A(_06895_),
    .X(_01244_));
 sky130_fd_sc_hd__mux2_1 _13644_ (.A0(\regs[28][29] ),
    .A1(_06353_),
    .S(_06886_),
    .X(_06896_));
 sky130_fd_sc_hd__clkbuf_1 _13645_ (.A(_06896_),
    .X(_01245_));
 sky130_fd_sc_hd__mux2_1 _13646_ (.A0(\regs[28][30] ),
    .A1(_06355_),
    .S(_06863_),
    .X(_06897_));
 sky130_fd_sc_hd__clkbuf_1 _13647_ (.A(_06897_),
    .X(_01246_));
 sky130_fd_sc_hd__mux2_1 _13648_ (.A0(\regs[28][31] ),
    .A1(_06357_),
    .S(_06863_),
    .X(_06898_));
 sky130_fd_sc_hd__clkbuf_1 _13649_ (.A(_06898_),
    .X(_01247_));
 sky130_fd_sc_hd__or2_4 _13650_ (.A(_04757_),
    .B(_05883_),
    .X(_06899_));
 sky130_fd_sc_hd__buf_6 _13651_ (.A(_06899_),
    .X(_06900_));
 sky130_fd_sc_hd__mux2_1 _13652_ (.A0(_05813_),
    .A1(\regs[2][0] ),
    .S(_06900_),
    .X(_06901_));
 sky130_fd_sc_hd__clkbuf_1 _13653_ (.A(_06901_),
    .X(_01248_));
 sky130_fd_sc_hd__mux2_1 _13654_ (.A0(_05819_),
    .A1(\regs[2][1] ),
    .S(_06900_),
    .X(_06902_));
 sky130_fd_sc_hd__clkbuf_1 _13655_ (.A(_06902_),
    .X(_01249_));
 sky130_fd_sc_hd__mux2_1 _13656_ (.A0(_05821_),
    .A1(\regs[2][2] ),
    .S(_06900_),
    .X(_06903_));
 sky130_fd_sc_hd__clkbuf_1 _13657_ (.A(_06903_),
    .X(_01250_));
 sky130_fd_sc_hd__mux2_1 _13658_ (.A0(_05823_),
    .A1(\regs[2][3] ),
    .S(_06900_),
    .X(_06904_));
 sky130_fd_sc_hd__clkbuf_1 _13659_ (.A(_06904_),
    .X(_01251_));
 sky130_fd_sc_hd__mux2_1 _13660_ (.A0(_05825_),
    .A1(\regs[2][4] ),
    .S(_06900_),
    .X(_06905_));
 sky130_fd_sc_hd__clkbuf_1 _13661_ (.A(_06905_),
    .X(_01252_));
 sky130_fd_sc_hd__mux2_1 _13662_ (.A0(_05827_),
    .A1(\regs[2][5] ),
    .S(_06900_),
    .X(_06906_));
 sky130_fd_sc_hd__clkbuf_1 _13663_ (.A(_06906_),
    .X(_01253_));
 sky130_fd_sc_hd__mux2_1 _13664_ (.A0(_05829_),
    .A1(\regs[2][6] ),
    .S(_06900_),
    .X(_06907_));
 sky130_fd_sc_hd__clkbuf_1 _13665_ (.A(_06907_),
    .X(_01254_));
 sky130_fd_sc_hd__mux2_1 _13666_ (.A0(_05831_),
    .A1(\regs[2][7] ),
    .S(_06900_),
    .X(_06908_));
 sky130_fd_sc_hd__clkbuf_1 _13667_ (.A(_06908_),
    .X(_01255_));
 sky130_fd_sc_hd__mux2_1 _13668_ (.A0(_05833_),
    .A1(\regs[2][8] ),
    .S(_06900_),
    .X(_06909_));
 sky130_fd_sc_hd__clkbuf_1 _13669_ (.A(_06909_),
    .X(_01256_));
 sky130_fd_sc_hd__mux2_1 _13670_ (.A0(_05835_),
    .A1(\regs[2][9] ),
    .S(_06900_),
    .X(_06910_));
 sky130_fd_sc_hd__clkbuf_1 _13671_ (.A(_06910_),
    .X(_01257_));
 sky130_fd_sc_hd__buf_6 _13672_ (.A(_06899_),
    .X(_06911_));
 sky130_fd_sc_hd__mux2_1 _13673_ (.A0(_05837_),
    .A1(\regs[2][10] ),
    .S(_06911_),
    .X(_06912_));
 sky130_fd_sc_hd__clkbuf_1 _13674_ (.A(_06912_),
    .X(_01258_));
 sky130_fd_sc_hd__mux2_1 _13675_ (.A0(_05840_),
    .A1(\regs[2][11] ),
    .S(_06911_),
    .X(_06913_));
 sky130_fd_sc_hd__clkbuf_1 _13676_ (.A(_06913_),
    .X(_01259_));
 sky130_fd_sc_hd__mux2_1 _13677_ (.A0(_05842_),
    .A1(\regs[2][12] ),
    .S(_06911_),
    .X(_06914_));
 sky130_fd_sc_hd__clkbuf_1 _13678_ (.A(_06914_),
    .X(_01260_));
 sky130_fd_sc_hd__mux2_1 _13679_ (.A0(_05844_),
    .A1(\regs[2][13] ),
    .S(_06911_),
    .X(_06915_));
 sky130_fd_sc_hd__clkbuf_1 _13680_ (.A(_06915_),
    .X(_01261_));
 sky130_fd_sc_hd__mux2_1 _13681_ (.A0(_05846_),
    .A1(\regs[2][14] ),
    .S(_06911_),
    .X(_06916_));
 sky130_fd_sc_hd__clkbuf_1 _13682_ (.A(_06916_),
    .X(_01262_));
 sky130_fd_sc_hd__mux2_1 _13683_ (.A0(_05848_),
    .A1(\regs[2][15] ),
    .S(_06911_),
    .X(_06917_));
 sky130_fd_sc_hd__clkbuf_1 _13684_ (.A(_06917_),
    .X(_01263_));
 sky130_fd_sc_hd__mux2_1 _13685_ (.A0(_05850_),
    .A1(\regs[2][16] ),
    .S(_06911_),
    .X(_06918_));
 sky130_fd_sc_hd__clkbuf_1 _13686_ (.A(_06918_),
    .X(_01264_));
 sky130_fd_sc_hd__mux2_1 _13687_ (.A0(_05852_),
    .A1(\regs[2][17] ),
    .S(_06911_),
    .X(_06919_));
 sky130_fd_sc_hd__clkbuf_1 _13688_ (.A(_06919_),
    .X(_01265_));
 sky130_fd_sc_hd__mux2_1 _13689_ (.A0(_05854_),
    .A1(\regs[2][18] ),
    .S(_06911_),
    .X(_06920_));
 sky130_fd_sc_hd__clkbuf_1 _13690_ (.A(_06920_),
    .X(_01266_));
 sky130_fd_sc_hd__mux2_1 _13691_ (.A0(_05856_),
    .A1(\regs[2][19] ),
    .S(_06911_),
    .X(_06921_));
 sky130_fd_sc_hd__clkbuf_1 _13692_ (.A(_06921_),
    .X(_01267_));
 sky130_fd_sc_hd__buf_6 _13693_ (.A(_06899_),
    .X(_06922_));
 sky130_fd_sc_hd__mux2_1 _13694_ (.A0(_05858_),
    .A1(\regs[2][20] ),
    .S(_06922_),
    .X(_06923_));
 sky130_fd_sc_hd__clkbuf_1 _13695_ (.A(_06923_),
    .X(_01268_));
 sky130_fd_sc_hd__mux2_1 _13696_ (.A0(_05861_),
    .A1(\regs[2][21] ),
    .S(_06922_),
    .X(_06924_));
 sky130_fd_sc_hd__clkbuf_1 _13697_ (.A(_06924_),
    .X(_01269_));
 sky130_fd_sc_hd__mux2_1 _13698_ (.A0(_05863_),
    .A1(\regs[2][22] ),
    .S(_06922_),
    .X(_06925_));
 sky130_fd_sc_hd__clkbuf_1 _13699_ (.A(_06925_),
    .X(_01270_));
 sky130_fd_sc_hd__mux2_1 _13700_ (.A0(_05865_),
    .A1(\regs[2][23] ),
    .S(_06922_),
    .X(_06926_));
 sky130_fd_sc_hd__clkbuf_1 _13701_ (.A(_06926_),
    .X(_01271_));
 sky130_fd_sc_hd__mux2_1 _13702_ (.A0(_05867_),
    .A1(\regs[2][24] ),
    .S(_06922_),
    .X(_06927_));
 sky130_fd_sc_hd__clkbuf_1 _13703_ (.A(_06927_),
    .X(_01272_));
 sky130_fd_sc_hd__mux2_1 _13704_ (.A0(_05869_),
    .A1(\regs[2][25] ),
    .S(_06922_),
    .X(_06928_));
 sky130_fd_sc_hd__clkbuf_1 _13705_ (.A(_06928_),
    .X(_01273_));
 sky130_fd_sc_hd__mux2_1 _13706_ (.A0(_05871_),
    .A1(\regs[2][26] ),
    .S(_06922_),
    .X(_06929_));
 sky130_fd_sc_hd__clkbuf_1 _13707_ (.A(_06929_),
    .X(_01274_));
 sky130_fd_sc_hd__mux2_1 _13708_ (.A0(_05873_),
    .A1(\regs[2][27] ),
    .S(_06922_),
    .X(_06930_));
 sky130_fd_sc_hd__clkbuf_1 _13709_ (.A(_06930_),
    .X(_01275_));
 sky130_fd_sc_hd__mux2_1 _13710_ (.A0(_05875_),
    .A1(\regs[2][28] ),
    .S(_06922_),
    .X(_06931_));
 sky130_fd_sc_hd__clkbuf_1 _13711_ (.A(_06931_),
    .X(_01276_));
 sky130_fd_sc_hd__mux2_1 _13712_ (.A0(_05877_),
    .A1(\regs[2][29] ),
    .S(_06922_),
    .X(_06932_));
 sky130_fd_sc_hd__clkbuf_1 _13713_ (.A(_06932_),
    .X(_01277_));
 sky130_fd_sc_hd__mux2_1 _13714_ (.A0(_05879_),
    .A1(\regs[2][30] ),
    .S(_06899_),
    .X(_06933_));
 sky130_fd_sc_hd__clkbuf_1 _13715_ (.A(_06933_),
    .X(_01278_));
 sky130_fd_sc_hd__mux2_1 _13716_ (.A0(_05881_),
    .A1(\regs[2][31] ),
    .S(_06899_),
    .X(_06934_));
 sky130_fd_sc_hd__clkbuf_1 _13717_ (.A(_06934_),
    .X(_01279_));
 sky130_fd_sc_hd__nor2_2 _13718_ (.A(_05883_),
    .B(_06218_),
    .Y(_06935_));
 sky130_fd_sc_hd__clkbuf_8 _13719_ (.A(_06935_),
    .X(_06936_));
 sky130_fd_sc_hd__mux2_1 _13720_ (.A0(\regs[30][0] ),
    .A1(_06291_),
    .S(_06936_),
    .X(_06937_));
 sky130_fd_sc_hd__clkbuf_1 _13721_ (.A(_06937_),
    .X(_01280_));
 sky130_fd_sc_hd__mux2_1 _13722_ (.A0(\regs[30][1] ),
    .A1(_06295_),
    .S(_06936_),
    .X(_06938_));
 sky130_fd_sc_hd__clkbuf_1 _13723_ (.A(_06938_),
    .X(_01281_));
 sky130_fd_sc_hd__mux2_1 _13724_ (.A0(\regs[30][2] ),
    .A1(_06297_),
    .S(_06936_),
    .X(_06939_));
 sky130_fd_sc_hd__clkbuf_1 _13725_ (.A(_06939_),
    .X(_01282_));
 sky130_fd_sc_hd__mux2_1 _13726_ (.A0(\regs[30][3] ),
    .A1(_06299_),
    .S(_06936_),
    .X(_06940_));
 sky130_fd_sc_hd__clkbuf_1 _13727_ (.A(_06940_),
    .X(_01283_));
 sky130_fd_sc_hd__mux2_1 _13728_ (.A0(\regs[30][4] ),
    .A1(_06301_),
    .S(_06936_),
    .X(_06941_));
 sky130_fd_sc_hd__clkbuf_1 _13729_ (.A(_06941_),
    .X(_01284_));
 sky130_fd_sc_hd__mux2_1 _13730_ (.A0(\regs[30][5] ),
    .A1(_06303_),
    .S(_06936_),
    .X(_06942_));
 sky130_fd_sc_hd__clkbuf_1 _13731_ (.A(_06942_),
    .X(_01285_));
 sky130_fd_sc_hd__mux2_1 _13732_ (.A0(\regs[30][6] ),
    .A1(_06305_),
    .S(_06936_),
    .X(_06943_));
 sky130_fd_sc_hd__clkbuf_1 _13733_ (.A(_06943_),
    .X(_01286_));
 sky130_fd_sc_hd__mux2_1 _13734_ (.A0(\regs[30][7] ),
    .A1(_06307_),
    .S(_06936_),
    .X(_06944_));
 sky130_fd_sc_hd__clkbuf_1 _13735_ (.A(_06944_),
    .X(_01287_));
 sky130_fd_sc_hd__mux2_1 _13736_ (.A0(\regs[30][8] ),
    .A1(_06309_),
    .S(_06936_),
    .X(_06945_));
 sky130_fd_sc_hd__clkbuf_1 _13737_ (.A(_06945_),
    .X(_01288_));
 sky130_fd_sc_hd__mux2_1 _13738_ (.A0(\regs[30][9] ),
    .A1(_06311_),
    .S(_06936_),
    .X(_06946_));
 sky130_fd_sc_hd__clkbuf_1 _13739_ (.A(_06946_),
    .X(_01289_));
 sky130_fd_sc_hd__buf_4 _13740_ (.A(_06935_),
    .X(_06947_));
 sky130_fd_sc_hd__mux2_1 _13741_ (.A0(\regs[30][10] ),
    .A1(_06313_),
    .S(_06947_),
    .X(_06948_));
 sky130_fd_sc_hd__clkbuf_1 _13742_ (.A(_06948_),
    .X(_01290_));
 sky130_fd_sc_hd__mux2_1 _13743_ (.A0(\regs[30][11] ),
    .A1(_06316_),
    .S(_06947_),
    .X(_06949_));
 sky130_fd_sc_hd__clkbuf_1 _13744_ (.A(_06949_),
    .X(_01291_));
 sky130_fd_sc_hd__mux2_1 _13745_ (.A0(\regs[30][12] ),
    .A1(_06318_),
    .S(_06947_),
    .X(_06950_));
 sky130_fd_sc_hd__clkbuf_1 _13746_ (.A(_06950_),
    .X(_01292_));
 sky130_fd_sc_hd__mux2_1 _13747_ (.A0(\regs[30][13] ),
    .A1(_06320_),
    .S(_06947_),
    .X(_06951_));
 sky130_fd_sc_hd__clkbuf_1 _13748_ (.A(_06951_),
    .X(_01293_));
 sky130_fd_sc_hd__mux2_1 _13749_ (.A0(\regs[30][14] ),
    .A1(_06322_),
    .S(_06947_),
    .X(_06952_));
 sky130_fd_sc_hd__clkbuf_1 _13750_ (.A(_06952_),
    .X(_01294_));
 sky130_fd_sc_hd__mux2_1 _13751_ (.A0(\regs[30][15] ),
    .A1(_06324_),
    .S(_06947_),
    .X(_06953_));
 sky130_fd_sc_hd__clkbuf_1 _13752_ (.A(_06953_),
    .X(_01295_));
 sky130_fd_sc_hd__mux2_1 _13753_ (.A0(\regs[30][16] ),
    .A1(_06326_),
    .S(_06947_),
    .X(_06954_));
 sky130_fd_sc_hd__clkbuf_1 _13754_ (.A(_06954_),
    .X(_01296_));
 sky130_fd_sc_hd__mux2_1 _13755_ (.A0(\regs[30][17] ),
    .A1(_06328_),
    .S(_06947_),
    .X(_06955_));
 sky130_fd_sc_hd__clkbuf_1 _13756_ (.A(_06955_),
    .X(_01297_));
 sky130_fd_sc_hd__mux2_1 _13757_ (.A0(\regs[30][18] ),
    .A1(_06330_),
    .S(_06947_),
    .X(_06956_));
 sky130_fd_sc_hd__clkbuf_1 _13758_ (.A(_06956_),
    .X(_01298_));
 sky130_fd_sc_hd__mux2_1 _13759_ (.A0(\regs[30][19] ),
    .A1(_06332_),
    .S(_06947_),
    .X(_06957_));
 sky130_fd_sc_hd__clkbuf_1 _13760_ (.A(_06957_),
    .X(_01299_));
 sky130_fd_sc_hd__buf_4 _13761_ (.A(_06935_),
    .X(_06958_));
 sky130_fd_sc_hd__mux2_1 _13762_ (.A0(\regs[30][20] ),
    .A1(_06334_),
    .S(_06958_),
    .X(_06959_));
 sky130_fd_sc_hd__clkbuf_1 _13763_ (.A(_06959_),
    .X(_01300_));
 sky130_fd_sc_hd__mux2_1 _13764_ (.A0(\regs[30][21] ),
    .A1(_06337_),
    .S(_06958_),
    .X(_06960_));
 sky130_fd_sc_hd__clkbuf_1 _13765_ (.A(_06960_),
    .X(_01301_));
 sky130_fd_sc_hd__mux2_1 _13766_ (.A0(\regs[30][22] ),
    .A1(_06339_),
    .S(_06958_),
    .X(_06961_));
 sky130_fd_sc_hd__clkbuf_1 _13767_ (.A(_06961_),
    .X(_01302_));
 sky130_fd_sc_hd__mux2_1 _13768_ (.A0(\regs[30][23] ),
    .A1(_06341_),
    .S(_06958_),
    .X(_06962_));
 sky130_fd_sc_hd__clkbuf_1 _13769_ (.A(_06962_),
    .X(_01303_));
 sky130_fd_sc_hd__mux2_1 _13770_ (.A0(\regs[30][24] ),
    .A1(_06343_),
    .S(_06958_),
    .X(_06963_));
 sky130_fd_sc_hd__clkbuf_1 _13771_ (.A(_06963_),
    .X(_01304_));
 sky130_fd_sc_hd__mux2_1 _13772_ (.A0(\regs[30][25] ),
    .A1(_06345_),
    .S(_06958_),
    .X(_06964_));
 sky130_fd_sc_hd__clkbuf_1 _13773_ (.A(_06964_),
    .X(_01305_));
 sky130_fd_sc_hd__mux2_1 _13774_ (.A0(\regs[30][26] ),
    .A1(_06347_),
    .S(_06958_),
    .X(_06965_));
 sky130_fd_sc_hd__clkbuf_1 _13775_ (.A(_06965_),
    .X(_01306_));
 sky130_fd_sc_hd__mux2_1 _13776_ (.A0(\regs[30][27] ),
    .A1(_06349_),
    .S(_06958_),
    .X(_06966_));
 sky130_fd_sc_hd__clkbuf_1 _13777_ (.A(_06966_),
    .X(_01307_));
 sky130_fd_sc_hd__mux2_1 _13778_ (.A0(\regs[30][28] ),
    .A1(_06351_),
    .S(_06958_),
    .X(_06967_));
 sky130_fd_sc_hd__clkbuf_1 _13779_ (.A(_06967_),
    .X(_01308_));
 sky130_fd_sc_hd__mux2_1 _13780_ (.A0(\regs[30][29] ),
    .A1(_06353_),
    .S(_06958_),
    .X(_06968_));
 sky130_fd_sc_hd__clkbuf_1 _13781_ (.A(_06968_),
    .X(_01309_));
 sky130_fd_sc_hd__mux2_1 _13782_ (.A0(\regs[30][30] ),
    .A1(_06355_),
    .S(_06935_),
    .X(_06969_));
 sky130_fd_sc_hd__clkbuf_1 _13783_ (.A(_06969_),
    .X(_01310_));
 sky130_fd_sc_hd__mux2_1 _13784_ (.A0(\regs[30][31] ),
    .A1(_06357_),
    .S(_06935_),
    .X(_06970_));
 sky130_fd_sc_hd__clkbuf_1 _13785_ (.A(_06970_),
    .X(_01311_));
 sky130_fd_sc_hd__inv_2 _13786_ (.A(_06070_),
    .Y(_00073_));
 sky130_fd_sc_hd__inv_2 _13787_ (.A(_06070_),
    .Y(_00074_));
 sky130_fd_sc_hd__inv_2 _13788_ (.A(_06070_),
    .Y(_00075_));
 sky130_fd_sc_hd__inv_2 _13789_ (.A(_06070_),
    .Y(_00076_));
 sky130_fd_sc_hd__inv_2 _13790_ (.A(_06070_),
    .Y(_00077_));
 sky130_fd_sc_hd__inv_2 _13791_ (.A(_06070_),
    .Y(_00078_));
 sky130_fd_sc_hd__buf_8 _13792_ (.A(_06069_),
    .X(_06971_));
 sky130_fd_sc_hd__inv_2 _13793_ (.A(_06971_),
    .Y(_00079_));
 sky130_fd_sc_hd__inv_2 _13794_ (.A(_06971_),
    .Y(_00080_));
 sky130_fd_sc_hd__inv_2 _13795_ (.A(_06971_),
    .Y(_00081_));
 sky130_fd_sc_hd__inv_2 _13796_ (.A(_06971_),
    .Y(_00082_));
 sky130_fd_sc_hd__inv_2 _13797_ (.A(_06971_),
    .Y(_00083_));
 sky130_fd_sc_hd__inv_2 _13798_ (.A(_06971_),
    .Y(_00084_));
 sky130_fd_sc_hd__inv_2 _13799_ (.A(_06971_),
    .Y(_00085_));
 sky130_fd_sc_hd__inv_2 _13800_ (.A(_06971_),
    .Y(_00086_));
 sky130_fd_sc_hd__inv_2 _13801_ (.A(_06971_),
    .Y(_00087_));
 sky130_fd_sc_hd__inv_2 _13802_ (.A(_06971_),
    .Y(_00088_));
 sky130_fd_sc_hd__buf_6 _13803_ (.A(_06069_),
    .X(_06972_));
 sky130_fd_sc_hd__inv_2 _13804_ (.A(_06972_),
    .Y(_00089_));
 sky130_fd_sc_hd__inv_2 _13805_ (.A(_06972_),
    .Y(_00090_));
 sky130_fd_sc_hd__inv_2 _13806_ (.A(_06972_),
    .Y(_00091_));
 sky130_fd_sc_hd__inv_2 _13807_ (.A(_06972_),
    .Y(_00092_));
 sky130_fd_sc_hd__inv_2 _13808_ (.A(_06972_),
    .Y(_00093_));
 sky130_fd_sc_hd__inv_2 _13809_ (.A(_06972_),
    .Y(_00094_));
 sky130_fd_sc_hd__inv_2 _13810_ (.A(_06972_),
    .Y(_00095_));
 sky130_fd_sc_hd__inv_2 _13811_ (.A(_06972_),
    .Y(_00096_));
 sky130_fd_sc_hd__inv_2 _13812_ (.A(_06972_),
    .Y(_00097_));
 sky130_fd_sc_hd__inv_2 _13813_ (.A(_06972_),
    .Y(_00098_));
 sky130_fd_sc_hd__buf_6 _13814_ (.A(_06069_),
    .X(_06973_));
 sky130_fd_sc_hd__inv_2 _13815_ (.A(_06973_),
    .Y(_00099_));
 sky130_fd_sc_hd__inv_2 _13816_ (.A(_06973_),
    .Y(_00100_));
 sky130_fd_sc_hd__inv_2 _13817_ (.A(_06973_),
    .Y(_00101_));
 sky130_fd_sc_hd__inv_2 _13818_ (.A(_06973_),
    .Y(_00102_));
 sky130_fd_sc_hd__inv_2 _13819_ (.A(_06973_),
    .Y(_00103_));
 sky130_fd_sc_hd__inv_2 _13820_ (.A(_06973_),
    .Y(_00104_));
 sky130_fd_sc_hd__inv_2 _13821_ (.A(_06973_),
    .Y(_00105_));
 sky130_fd_sc_hd__inv_2 _13822_ (.A(_06973_),
    .Y(_00106_));
 sky130_fd_sc_hd__inv_2 _13823_ (.A(_06973_),
    .Y(_00107_));
 sky130_fd_sc_hd__inv_2 _13824_ (.A(_06973_),
    .Y(_00108_));
 sky130_fd_sc_hd__buf_4 _13825_ (.A(_06069_),
    .X(_06974_));
 sky130_fd_sc_hd__inv_2 _13826_ (.A(_06974_),
    .Y(_00109_));
 sky130_fd_sc_hd__inv_2 _13827_ (.A(_06974_),
    .Y(_00110_));
 sky130_fd_sc_hd__inv_2 _13828_ (.A(_06974_),
    .Y(_00111_));
 sky130_fd_sc_hd__inv_2 _13829_ (.A(_06974_),
    .Y(_00112_));
 sky130_fd_sc_hd__inv_2 _13830_ (.A(_06974_),
    .Y(_00113_));
 sky130_fd_sc_hd__inv_2 _13831_ (.A(_06974_),
    .Y(_00114_));
 sky130_fd_sc_hd__inv_2 _13832_ (.A(_06974_),
    .Y(_00115_));
 sky130_fd_sc_hd__inv_2 _13833_ (.A(_06974_),
    .Y(_00116_));
 sky130_fd_sc_hd__inv_2 _13834_ (.A(_06974_),
    .Y(_00117_));
 sky130_fd_sc_hd__inv_2 _13835_ (.A(_06974_),
    .Y(_00118_));
 sky130_fd_sc_hd__buf_4 _13836_ (.A(_06069_),
    .X(_06975_));
 sky130_fd_sc_hd__inv_2 _13837_ (.A(_06975_),
    .Y(_00119_));
 sky130_fd_sc_hd__inv_2 _13838_ (.A(_06975_),
    .Y(_00120_));
 sky130_fd_sc_hd__inv_2 _13839_ (.A(_06975_),
    .Y(_00121_));
 sky130_fd_sc_hd__inv_2 _13840_ (.A(_06975_),
    .Y(_00122_));
 sky130_fd_sc_hd__inv_2 _13841_ (.A(_06975_),
    .Y(_00123_));
 sky130_fd_sc_hd__inv_2 _13842_ (.A(_06975_),
    .Y(_00124_));
 sky130_fd_sc_hd__inv_2 _13843_ (.A(_06975_),
    .Y(_00125_));
 sky130_fd_sc_hd__inv_2 _13844_ (.A(_06975_),
    .Y(_00126_));
 sky130_fd_sc_hd__inv_2 _13845_ (.A(_06975_),
    .Y(_00127_));
 sky130_fd_sc_hd__inv_2 _13846_ (.A(_06975_),
    .Y(_00128_));
 sky130_fd_sc_hd__buf_4 _13847_ (.A(_06069_),
    .X(_06976_));
 sky130_fd_sc_hd__inv_2 _13848_ (.A(_06976_),
    .Y(_00129_));
 sky130_fd_sc_hd__inv_2 _13849_ (.A(_06976_),
    .Y(_00130_));
 sky130_fd_sc_hd__inv_2 _13850_ (.A(_06976_),
    .Y(_00131_));
 sky130_fd_sc_hd__inv_2 _13851_ (.A(_06976_),
    .Y(_00132_));
 sky130_fd_sc_hd__inv_2 _13852_ (.A(_06976_),
    .Y(_00133_));
 sky130_fd_sc_hd__inv_2 _13853_ (.A(_06976_),
    .Y(_00134_));
 sky130_fd_sc_hd__inv_2 _13854_ (.A(_06976_),
    .Y(_00135_));
 sky130_fd_sc_hd__inv_2 _13855_ (.A(_06976_),
    .Y(_00136_));
 sky130_fd_sc_hd__inv_2 _13856_ (.A(_06976_),
    .Y(_00137_));
 sky130_fd_sc_hd__inv_2 _13857_ (.A(_06976_),
    .Y(_00138_));
 sky130_fd_sc_hd__buf_4 _13858_ (.A(_06069_),
    .X(_06977_));
 sky130_fd_sc_hd__inv_2 _13859_ (.A(_06977_),
    .Y(_00139_));
 sky130_fd_sc_hd__inv_2 _13860_ (.A(_06977_),
    .Y(_00140_));
 sky130_fd_sc_hd__inv_2 _13861_ (.A(_06977_),
    .Y(_00141_));
 sky130_fd_sc_hd__inv_2 _13862_ (.A(_06977_),
    .Y(_00142_));
 sky130_fd_sc_hd__inv_2 _13863_ (.A(_06977_),
    .Y(_00143_));
 sky130_fd_sc_hd__inv_2 _13864_ (.A(_06977_),
    .Y(_00144_));
 sky130_fd_sc_hd__inv_2 _13865_ (.A(_06977_),
    .Y(_00145_));
 sky130_fd_sc_hd__inv_2 _13866_ (.A(_06977_),
    .Y(_00146_));
 sky130_fd_sc_hd__inv_2 _13867_ (.A(_06977_),
    .Y(_00147_));
 sky130_fd_sc_hd__inv_2 _13868_ (.A(_06977_),
    .Y(_00148_));
 sky130_fd_sc_hd__buf_4 _13869_ (.A(_06069_),
    .X(_06978_));
 sky130_fd_sc_hd__inv_2 _13870_ (.A(_06978_),
    .Y(_00149_));
 sky130_fd_sc_hd__inv_2 _13871_ (.A(_06978_),
    .Y(_00150_));
 sky130_fd_sc_hd__inv_2 _13872_ (.A(_06978_),
    .Y(_00151_));
 sky130_fd_sc_hd__inv_2 _13873_ (.A(_06978_),
    .Y(_00152_));
 sky130_fd_sc_hd__inv_2 _13874_ (.A(_06978_),
    .Y(_00153_));
 sky130_fd_sc_hd__inv_2 _13875_ (.A(_06978_),
    .Y(_00154_));
 sky130_fd_sc_hd__inv_2 _13876_ (.A(_06978_),
    .Y(_00155_));
 sky130_fd_sc_hd__inv_2 _13877_ (.A(_06978_),
    .Y(_00156_));
 sky130_fd_sc_hd__inv_2 _13878_ (.A(_06978_),
    .Y(_00157_));
 sky130_fd_sc_hd__inv_2 _13879_ (.A(_06978_),
    .Y(_00158_));
 sky130_fd_sc_hd__buf_4 _13880_ (.A(_06069_),
    .X(_06979_));
 sky130_fd_sc_hd__inv_2 _13881_ (.A(_06979_),
    .Y(_00159_));
 sky130_fd_sc_hd__inv_2 _13882_ (.A(_06979_),
    .Y(_00160_));
 sky130_fd_sc_hd__inv_2 _13883_ (.A(_06979_),
    .Y(_00161_));
 sky130_fd_sc_hd__inv_2 _13884_ (.A(_06979_),
    .Y(_00162_));
 sky130_fd_sc_hd__inv_2 _13885_ (.A(_06979_),
    .Y(_00163_));
 sky130_fd_sc_hd__inv_2 _13886_ (.A(_06979_),
    .Y(_00164_));
 sky130_fd_sc_hd__inv_2 _13887_ (.A(_06979_),
    .Y(_00165_));
 sky130_fd_sc_hd__inv_2 _13888_ (.A(_06979_),
    .Y(_00166_));
 sky130_fd_sc_hd__inv_2 _13889_ (.A(_06979_),
    .Y(_00167_));
 sky130_fd_sc_hd__inv_2 _13890_ (.A(_06979_),
    .Y(_00168_));
 sky130_fd_sc_hd__buf_4 _13891_ (.A(_04755_),
    .X(_06980_));
 sky130_fd_sc_hd__clkbuf_8 _13892_ (.A(_06980_),
    .X(_06981_));
 sky130_fd_sc_hd__inv_2 _13893_ (.A(_06981_),
    .Y(_00169_));
 sky130_fd_sc_hd__inv_2 _13894_ (.A(_06981_),
    .Y(_00170_));
 sky130_fd_sc_hd__inv_2 _13895_ (.A(_06981_),
    .Y(_00171_));
 sky130_fd_sc_hd__inv_2 _13896_ (.A(_06981_),
    .Y(_00172_));
 sky130_fd_sc_hd__inv_2 _13897_ (.A(_06981_),
    .Y(_00173_));
 sky130_fd_sc_hd__inv_2 _13898_ (.A(_06981_),
    .Y(_00174_));
 sky130_fd_sc_hd__inv_2 _13899_ (.A(_06981_),
    .Y(_00175_));
 sky130_fd_sc_hd__inv_2 _13900_ (.A(_06981_),
    .Y(_00176_));
 sky130_fd_sc_hd__inv_2 _13901_ (.A(_06981_),
    .Y(_00177_));
 sky130_fd_sc_hd__inv_2 _13902_ (.A(_06981_),
    .Y(_00178_));
 sky130_fd_sc_hd__buf_4 _13903_ (.A(_06980_),
    .X(_06982_));
 sky130_fd_sc_hd__inv_2 _13904_ (.A(_06982_),
    .Y(_00179_));
 sky130_fd_sc_hd__inv_2 _13905_ (.A(_06982_),
    .Y(_00180_));
 sky130_fd_sc_hd__inv_2 _13906_ (.A(_06982_),
    .Y(_00181_));
 sky130_fd_sc_hd__inv_2 _13907_ (.A(_06982_),
    .Y(_00182_));
 sky130_fd_sc_hd__inv_2 _13908_ (.A(_06982_),
    .Y(_00183_));
 sky130_fd_sc_hd__inv_2 _13909_ (.A(_06982_),
    .Y(_00184_));
 sky130_fd_sc_hd__inv_2 _13910_ (.A(_06982_),
    .Y(_00185_));
 sky130_fd_sc_hd__inv_2 _13911_ (.A(_06982_),
    .Y(_00186_));
 sky130_fd_sc_hd__inv_2 _13912_ (.A(_06982_),
    .Y(_00187_));
 sky130_fd_sc_hd__inv_2 _13913_ (.A(_06982_),
    .Y(_00188_));
 sky130_fd_sc_hd__buf_4 _13914_ (.A(_06980_),
    .X(_06983_));
 sky130_fd_sc_hd__inv_2 _13915_ (.A(_06983_),
    .Y(_00189_));
 sky130_fd_sc_hd__inv_2 _13916_ (.A(_06983_),
    .Y(_00190_));
 sky130_fd_sc_hd__inv_2 _13917_ (.A(_06983_),
    .Y(_00191_));
 sky130_fd_sc_hd__inv_2 _13918_ (.A(_06983_),
    .Y(_00192_));
 sky130_fd_sc_hd__inv_2 _13919_ (.A(_06983_),
    .Y(_00193_));
 sky130_fd_sc_hd__inv_2 _13920_ (.A(_06983_),
    .Y(_00194_));
 sky130_fd_sc_hd__inv_2 _13921_ (.A(_06983_),
    .Y(_00195_));
 sky130_fd_sc_hd__inv_2 _13922_ (.A(_06983_),
    .Y(_00196_));
 sky130_fd_sc_hd__inv_2 _13923_ (.A(_06983_),
    .Y(_00197_));
 sky130_fd_sc_hd__inv_2 _13924_ (.A(_06983_),
    .Y(_00198_));
 sky130_fd_sc_hd__buf_6 _13925_ (.A(_06980_),
    .X(_06984_));
 sky130_fd_sc_hd__inv_2 _13926_ (.A(_06984_),
    .Y(_00199_));
 sky130_fd_sc_hd__inv_2 _13927_ (.A(_06984_),
    .Y(_00200_));
 sky130_fd_sc_hd__inv_2 _13928_ (.A(_06984_),
    .Y(_00201_));
 sky130_fd_sc_hd__inv_2 _13929_ (.A(_06984_),
    .Y(_00202_));
 sky130_fd_sc_hd__inv_2 _13930_ (.A(_06984_),
    .Y(_00203_));
 sky130_fd_sc_hd__inv_2 _13931_ (.A(_06984_),
    .Y(_00204_));
 sky130_fd_sc_hd__inv_2 _13932_ (.A(_06984_),
    .Y(_00205_));
 sky130_fd_sc_hd__inv_2 _13933_ (.A(_06984_),
    .Y(_00206_));
 sky130_fd_sc_hd__inv_2 _13934_ (.A(_06984_),
    .Y(_00207_));
 sky130_fd_sc_hd__inv_2 _13935_ (.A(_06984_),
    .Y(_00208_));
 sky130_fd_sc_hd__buf_4 _13936_ (.A(_06980_),
    .X(_06985_));
 sky130_fd_sc_hd__inv_2 _13937_ (.A(_06985_),
    .Y(_00209_));
 sky130_fd_sc_hd__inv_2 _13938_ (.A(_06985_),
    .Y(_00210_));
 sky130_fd_sc_hd__inv_2 _13939_ (.A(_06985_),
    .Y(_00211_));
 sky130_fd_sc_hd__inv_2 _13940_ (.A(_06985_),
    .Y(_00212_));
 sky130_fd_sc_hd__inv_2 _13941_ (.A(_06985_),
    .Y(_00213_));
 sky130_fd_sc_hd__inv_2 _13942_ (.A(_06985_),
    .Y(_00214_));
 sky130_fd_sc_hd__inv_2 _13943_ (.A(_06985_),
    .Y(_00215_));
 sky130_fd_sc_hd__inv_2 _13944_ (.A(_06985_),
    .Y(_00216_));
 sky130_fd_sc_hd__inv_2 _13945_ (.A(_06985_),
    .Y(_00217_));
 sky130_fd_sc_hd__inv_2 _13946_ (.A(_06985_),
    .Y(_00218_));
 sky130_fd_sc_hd__buf_4 _13947_ (.A(_06980_),
    .X(_06986_));
 sky130_fd_sc_hd__inv_2 _13948_ (.A(_06986_),
    .Y(_00219_));
 sky130_fd_sc_hd__inv_2 _13949_ (.A(_06986_),
    .Y(_00220_));
 sky130_fd_sc_hd__inv_2 _13950_ (.A(_06986_),
    .Y(_00221_));
 sky130_fd_sc_hd__inv_2 _13951_ (.A(_06986_),
    .Y(_00222_));
 sky130_fd_sc_hd__inv_2 _13952_ (.A(_06986_),
    .Y(_00223_));
 sky130_fd_sc_hd__inv_2 _13953_ (.A(_06986_),
    .Y(_00224_));
 sky130_fd_sc_hd__inv_2 _13954_ (.A(_06986_),
    .Y(_00225_));
 sky130_fd_sc_hd__inv_2 _13955_ (.A(_06986_),
    .Y(_00226_));
 sky130_fd_sc_hd__inv_2 _13956_ (.A(_06986_),
    .Y(_00227_));
 sky130_fd_sc_hd__inv_2 _13957_ (.A(_06986_),
    .Y(_00228_));
 sky130_fd_sc_hd__buf_4 _13958_ (.A(_06980_),
    .X(_06987_));
 sky130_fd_sc_hd__inv_2 _13959_ (.A(_06987_),
    .Y(_00229_));
 sky130_fd_sc_hd__inv_2 _13960_ (.A(_06987_),
    .Y(_00230_));
 sky130_fd_sc_hd__inv_2 _13961_ (.A(_06987_),
    .Y(_00231_));
 sky130_fd_sc_hd__inv_2 _13962_ (.A(_06987_),
    .Y(_00232_));
 sky130_fd_sc_hd__inv_2 _13963_ (.A(_06987_),
    .Y(_00233_));
 sky130_fd_sc_hd__inv_2 _13964_ (.A(_06987_),
    .Y(_00234_));
 sky130_fd_sc_hd__inv_2 _13965_ (.A(_06987_),
    .Y(_00235_));
 sky130_fd_sc_hd__inv_2 _13966_ (.A(_06987_),
    .Y(_00236_));
 sky130_fd_sc_hd__inv_2 _13967_ (.A(_06987_),
    .Y(_00237_));
 sky130_fd_sc_hd__inv_2 _13968_ (.A(_06987_),
    .Y(_00238_));
 sky130_fd_sc_hd__buf_4 _13969_ (.A(_06980_),
    .X(_06988_));
 sky130_fd_sc_hd__inv_2 _13970_ (.A(_06988_),
    .Y(_00239_));
 sky130_fd_sc_hd__inv_2 _13971_ (.A(_06988_),
    .Y(_00240_));
 sky130_fd_sc_hd__inv_2 _13972_ (.A(_06988_),
    .Y(_00241_));
 sky130_fd_sc_hd__inv_2 _13973_ (.A(_06988_),
    .Y(_00242_));
 sky130_fd_sc_hd__inv_2 _13974_ (.A(_06988_),
    .Y(_00243_));
 sky130_fd_sc_hd__inv_2 _13975_ (.A(_06988_),
    .Y(_00244_));
 sky130_fd_sc_hd__inv_2 _13976_ (.A(_06988_),
    .Y(_00245_));
 sky130_fd_sc_hd__inv_2 _13977_ (.A(_06988_),
    .Y(_00246_));
 sky130_fd_sc_hd__inv_2 _13978_ (.A(_06988_),
    .Y(_00247_));
 sky130_fd_sc_hd__inv_2 _13979_ (.A(_06988_),
    .Y(_00248_));
 sky130_fd_sc_hd__buf_4 _13980_ (.A(_06980_),
    .X(_06989_));
 sky130_fd_sc_hd__inv_2 _13981_ (.A(_06989_),
    .Y(_00249_));
 sky130_fd_sc_hd__inv_2 _13982_ (.A(_06989_),
    .Y(_00250_));
 sky130_fd_sc_hd__inv_2 _13983_ (.A(_06989_),
    .Y(_00251_));
 sky130_fd_sc_hd__inv_2 _13984_ (.A(_06989_),
    .Y(_00252_));
 sky130_fd_sc_hd__inv_2 _13985_ (.A(_06989_),
    .Y(_00253_));
 sky130_fd_sc_hd__inv_2 _13986_ (.A(_06989_),
    .Y(_00254_));
 sky130_fd_sc_hd__inv_2 _13987_ (.A(_06989_),
    .Y(_00255_));
 sky130_fd_sc_hd__inv_2 _13988_ (.A(_06989_),
    .Y(_00256_));
 sky130_fd_sc_hd__inv_2 _13989_ (.A(_06989_),
    .Y(_00257_));
 sky130_fd_sc_hd__inv_2 _13990_ (.A(_06989_),
    .Y(_00258_));
 sky130_fd_sc_hd__buf_4 _13991_ (.A(_06980_),
    .X(_06990_));
 sky130_fd_sc_hd__inv_2 _13992_ (.A(_06990_),
    .Y(_00259_));
 sky130_fd_sc_hd__inv_2 _13993_ (.A(_06990_),
    .Y(_00260_));
 sky130_fd_sc_hd__inv_2 _13994_ (.A(_06990_),
    .Y(_00261_));
 sky130_fd_sc_hd__inv_2 _13995_ (.A(_06990_),
    .Y(_00262_));
 sky130_fd_sc_hd__inv_2 _13996_ (.A(_06990_),
    .Y(_00263_));
 sky130_fd_sc_hd__inv_2 _13997_ (.A(_06990_),
    .Y(_00264_));
 sky130_fd_sc_hd__inv_2 _13998_ (.A(_06990_),
    .Y(_00265_));
 sky130_fd_sc_hd__inv_2 _13999_ (.A(_06990_),
    .Y(_00266_));
 sky130_fd_sc_hd__inv_2 _14000_ (.A(_06990_),
    .Y(_00267_));
 sky130_fd_sc_hd__inv_2 _14001_ (.A(_06990_),
    .Y(_00268_));
 sky130_fd_sc_hd__buf_4 _14002_ (.A(_04755_),
    .X(_06991_));
 sky130_fd_sc_hd__inv_2 _14003_ (.A(_06991_),
    .Y(_00269_));
 sky130_fd_sc_hd__inv_2 _14004_ (.A(_06991_),
    .Y(_00270_));
 sky130_fd_sc_hd__inv_2 _14005_ (.A(_06991_),
    .Y(_00271_));
 sky130_fd_sc_hd__inv_2 _14006_ (.A(_06991_),
    .Y(_00272_));
 sky130_fd_sc_hd__inv_2 _14007_ (.A(_06991_),
    .Y(_00273_));
 sky130_fd_sc_hd__inv_2 _14008_ (.A(_06991_),
    .Y(_00274_));
 sky130_fd_sc_hd__inv_2 _14009_ (.A(_06991_),
    .Y(_00275_));
 sky130_fd_sc_hd__inv_2 _14010_ (.A(_06991_),
    .Y(_00276_));
 sky130_fd_sc_hd__inv_2 _14011_ (.A(_06991_),
    .Y(_00277_));
 sky130_fd_sc_hd__inv_2 _14012_ (.A(_06991_),
    .Y(_00278_));
 sky130_fd_sc_hd__buf_4 _14013_ (.A(_04755_),
    .X(_06992_));
 sky130_fd_sc_hd__inv_2 _14014_ (.A(_06992_),
    .Y(_00279_));
 sky130_fd_sc_hd__inv_2 _14015_ (.A(_06992_),
    .Y(_00280_));
 sky130_fd_sc_hd__inv_2 _14016_ (.A(_06992_),
    .Y(_00281_));
 sky130_fd_sc_hd__inv_2 _14017_ (.A(_06992_),
    .Y(_00282_));
 sky130_fd_sc_hd__inv_2 _14018_ (.A(_06992_),
    .Y(_00283_));
 sky130_fd_sc_hd__inv_2 _14019_ (.A(_06992_),
    .Y(_00284_));
 sky130_fd_sc_hd__inv_2 _14020_ (.A(_06992_),
    .Y(_00285_));
 sky130_fd_sc_hd__inv_2 _14021_ (.A(_06992_),
    .Y(_00286_));
 sky130_fd_sc_hd__inv_2 _14022_ (.A(_06992_),
    .Y(_00287_));
 sky130_fd_sc_hd__inv_2 _14023_ (.A(_06992_),
    .Y(_00288_));
 sky130_fd_sc_hd__buf_4 _14024_ (.A(_04755_),
    .X(_06993_));
 sky130_fd_sc_hd__inv_2 _14025_ (.A(_06993_),
    .Y(_00289_));
 sky130_fd_sc_hd__inv_2 _14026_ (.A(_06993_),
    .Y(_00290_));
 sky130_fd_sc_hd__inv_2 _14027_ (.A(_06993_),
    .Y(_00291_));
 sky130_fd_sc_hd__inv_2 _14028_ (.A(_06993_),
    .Y(_00292_));
 sky130_fd_sc_hd__inv_2 _14029_ (.A(_06993_),
    .Y(_00293_));
 sky130_fd_sc_hd__inv_2 _14030_ (.A(_06993_),
    .Y(_00294_));
 sky130_fd_sc_hd__inv_2 _14031_ (.A(_06993_),
    .Y(_00295_));
 sky130_fd_sc_hd__inv_2 _14032_ (.A(_06993_),
    .Y(_00296_));
 sky130_fd_sc_hd__nor2_4 _14033_ (.A(_06072_),
    .B(_06145_),
    .Y(_06994_));
 sky130_fd_sc_hd__buf_6 _14034_ (.A(_06994_),
    .X(_06995_));
 sky130_fd_sc_hd__mux2_1 _14035_ (.A0(\regs[17][0] ),
    .A1(_04761_),
    .S(_06995_),
    .X(_06996_));
 sky130_fd_sc_hd__clkbuf_1 _14036_ (.A(_06996_),
    .X(_01472_));
 sky130_fd_sc_hd__mux2_1 _14037_ (.A0(\regs[17][1] ),
    .A1(_04817_),
    .S(_06995_),
    .X(_06997_));
 sky130_fd_sc_hd__clkbuf_1 _14038_ (.A(_06997_),
    .X(_01473_));
 sky130_fd_sc_hd__mux2_1 _14039_ (.A0(\regs[17][2] ),
    .A1(_04857_),
    .S(_06995_),
    .X(_06998_));
 sky130_fd_sc_hd__clkbuf_1 _14040_ (.A(_06998_),
    .X(_01474_));
 sky130_fd_sc_hd__mux2_1 _14041_ (.A0(\regs[17][3] ),
    .A1(_04903_),
    .S(_06995_),
    .X(_06999_));
 sky130_fd_sc_hd__clkbuf_1 _14042_ (.A(_06999_),
    .X(_01475_));
 sky130_fd_sc_hd__mux2_1 _14043_ (.A0(\regs[17][4] ),
    .A1(_04951_),
    .S(_06995_),
    .X(_07000_));
 sky130_fd_sc_hd__clkbuf_1 _14044_ (.A(_07000_),
    .X(_01476_));
 sky130_fd_sc_hd__mux2_1 _14045_ (.A0(\regs[17][5] ),
    .A1(_04991_),
    .S(_06995_),
    .X(_07001_));
 sky130_fd_sc_hd__clkbuf_1 _14046_ (.A(_07001_),
    .X(_01477_));
 sky130_fd_sc_hd__mux2_1 _14047_ (.A0(\regs[17][6] ),
    .A1(_05029_),
    .S(_06995_),
    .X(_07002_));
 sky130_fd_sc_hd__clkbuf_1 _14048_ (.A(_07002_),
    .X(_01478_));
 sky130_fd_sc_hd__mux2_1 _14049_ (.A0(\regs[17][7] ),
    .A1(_05079_),
    .S(_06995_),
    .X(_07003_));
 sky130_fd_sc_hd__clkbuf_1 _14050_ (.A(_07003_),
    .X(_01479_));
 sky130_fd_sc_hd__mux2_1 _14051_ (.A0(\regs[17][8] ),
    .A1(_05120_),
    .S(_06995_),
    .X(_07004_));
 sky130_fd_sc_hd__clkbuf_1 _14052_ (.A(_07004_),
    .X(_01480_));
 sky130_fd_sc_hd__mux2_1 _14053_ (.A0(\regs[17][9] ),
    .A1(_05156_),
    .S(_06995_),
    .X(_07005_));
 sky130_fd_sc_hd__clkbuf_1 _14054_ (.A(_07005_),
    .X(_01481_));
 sky130_fd_sc_hd__buf_6 _14055_ (.A(_06994_),
    .X(_07006_));
 sky130_fd_sc_hd__mux2_1 _14056_ (.A0(\regs[17][10] ),
    .A1(_05186_),
    .S(_07006_),
    .X(_07007_));
 sky130_fd_sc_hd__clkbuf_1 _14057_ (.A(_07007_),
    .X(_01482_));
 sky130_fd_sc_hd__mux2_1 _14058_ (.A0(\regs[17][11] ),
    .A1(_05223_),
    .S(_07006_),
    .X(_07008_));
 sky130_fd_sc_hd__clkbuf_1 _14059_ (.A(_07008_),
    .X(_01483_));
 sky130_fd_sc_hd__mux2_1 _14060_ (.A0(\regs[17][12] ),
    .A1(_05262_),
    .S(_07006_),
    .X(_07009_));
 sky130_fd_sc_hd__clkbuf_1 _14061_ (.A(_07009_),
    .X(_01484_));
 sky130_fd_sc_hd__mux2_1 _14062_ (.A0(\regs[17][13] ),
    .A1(_05295_),
    .S(_07006_),
    .X(_07010_));
 sky130_fd_sc_hd__clkbuf_1 _14063_ (.A(_07010_),
    .X(_01485_));
 sky130_fd_sc_hd__mux2_1 _14064_ (.A0(\regs[17][14] ),
    .A1(_05328_),
    .S(_07006_),
    .X(_07011_));
 sky130_fd_sc_hd__clkbuf_1 _14065_ (.A(_07011_),
    .X(_01486_));
 sky130_fd_sc_hd__mux2_1 _14066_ (.A0(\regs[17][15] ),
    .A1(_05358_),
    .S(_07006_),
    .X(_07012_));
 sky130_fd_sc_hd__clkbuf_1 _14067_ (.A(_07012_),
    .X(_01487_));
 sky130_fd_sc_hd__mux2_1 _14068_ (.A0(\regs[17][16] ),
    .A1(_05399_),
    .S(_07006_),
    .X(_07013_));
 sky130_fd_sc_hd__clkbuf_1 _14069_ (.A(_07013_),
    .X(_01488_));
 sky130_fd_sc_hd__mux2_1 _14070_ (.A0(\regs[17][17] ),
    .A1(_05423_),
    .S(_07006_),
    .X(_07014_));
 sky130_fd_sc_hd__clkbuf_1 _14071_ (.A(_07014_),
    .X(_01489_));
 sky130_fd_sc_hd__mux2_1 _14072_ (.A0(\regs[17][18] ),
    .A1(_05451_),
    .S(_07006_),
    .X(_07015_));
 sky130_fd_sc_hd__clkbuf_1 _14073_ (.A(_07015_),
    .X(_01490_));
 sky130_fd_sc_hd__mux2_1 _14074_ (.A0(\regs[17][19] ),
    .A1(_05476_),
    .S(_07006_),
    .X(_07016_));
 sky130_fd_sc_hd__clkbuf_1 _14075_ (.A(_07016_),
    .X(_01491_));
 sky130_fd_sc_hd__buf_4 _14076_ (.A(_06994_),
    .X(_07017_));
 sky130_fd_sc_hd__mux2_1 _14077_ (.A0(\regs[17][20] ),
    .A1(_05513_),
    .S(_07017_),
    .X(_07018_));
 sky130_fd_sc_hd__clkbuf_1 _14078_ (.A(_07018_),
    .X(_01492_));
 sky130_fd_sc_hd__mux2_1 _14079_ (.A0(\regs[17][21] ),
    .A1(_05540_),
    .S(_07017_),
    .X(_07019_));
 sky130_fd_sc_hd__clkbuf_1 _14080_ (.A(_07019_),
    .X(_01493_));
 sky130_fd_sc_hd__mux2_1 _14081_ (.A0(\regs[17][22] ),
    .A1(_05569_),
    .S(_07017_),
    .X(_07020_));
 sky130_fd_sc_hd__clkbuf_1 _14082_ (.A(_07020_),
    .X(_01494_));
 sky130_fd_sc_hd__mux2_1 _14083_ (.A0(\regs[17][23] ),
    .A1(_05599_),
    .S(_07017_),
    .X(_07021_));
 sky130_fd_sc_hd__clkbuf_1 _14084_ (.A(_07021_),
    .X(_01495_));
 sky130_fd_sc_hd__mux2_1 _14085_ (.A0(\regs[17][24] ),
    .A1(_05635_),
    .S(_07017_),
    .X(_07022_));
 sky130_fd_sc_hd__clkbuf_1 _14086_ (.A(_07022_),
    .X(_01496_));
 sky130_fd_sc_hd__mux2_1 _14087_ (.A0(\regs[17][25] ),
    .A1(_05659_),
    .S(_07017_),
    .X(_07023_));
 sky130_fd_sc_hd__clkbuf_1 _14088_ (.A(_07023_),
    .X(_01497_));
 sky130_fd_sc_hd__mux2_1 _14089_ (.A0(\regs[17][26] ),
    .A1(_05683_),
    .S(_07017_),
    .X(_07024_));
 sky130_fd_sc_hd__clkbuf_1 _14090_ (.A(_07024_),
    .X(_01498_));
 sky130_fd_sc_hd__mux2_1 _14091_ (.A0(\regs[17][27] ),
    .A1(_05707_),
    .S(_07017_),
    .X(_07025_));
 sky130_fd_sc_hd__clkbuf_1 _14092_ (.A(_07025_),
    .X(_01499_));
 sky130_fd_sc_hd__mux2_1 _14093_ (.A0(\regs[17][28] ),
    .A1(_05734_),
    .S(_07017_),
    .X(_07026_));
 sky130_fd_sc_hd__clkbuf_1 _14094_ (.A(_07026_),
    .X(_01500_));
 sky130_fd_sc_hd__mux2_1 _14095_ (.A0(\regs[17][29] ),
    .A1(_05762_),
    .S(_07017_),
    .X(_07027_));
 sky130_fd_sc_hd__clkbuf_1 _14096_ (.A(_07027_),
    .X(_01501_));
 sky130_fd_sc_hd__mux2_1 _14097_ (.A0(\regs[17][30] ),
    .A1(_05786_),
    .S(_06994_),
    .X(_07028_));
 sky130_fd_sc_hd__clkbuf_1 _14098_ (.A(_07028_),
    .X(_01502_));
 sky130_fd_sc_hd__mux2_1 _14099_ (.A0(\regs[17][31] ),
    .A1(_05810_),
    .S(_06994_),
    .X(_07029_));
 sky130_fd_sc_hd__clkbuf_1 _14100_ (.A(_07029_),
    .X(_01503_));
 sky130_fd_sc_hd__inv_2 _14101_ (.A(_06993_),
    .Y(_00297_));
 sky130_fd_sc_hd__inv_2 _14102_ (.A(_06993_),
    .Y(_00298_));
 sky130_fd_sc_hd__clkbuf_8 _14103_ (.A(_04755_),
    .X(_07030_));
 sky130_fd_sc_hd__inv_2 _14104_ (.A(_07030_),
    .Y(_00299_));
 sky130_fd_sc_hd__inv_2 _14105_ (.A(_07030_),
    .Y(_00300_));
 sky130_fd_sc_hd__inv_2 _14106_ (.A(_07030_),
    .Y(_00301_));
 sky130_fd_sc_hd__inv_2 _14107_ (.A(_07030_),
    .Y(_00302_));
 sky130_fd_sc_hd__inv_2 _14108_ (.A(_07030_),
    .Y(_00303_));
 sky130_fd_sc_hd__inv_2 _14109_ (.A(_07030_),
    .Y(_00304_));
 sky130_fd_sc_hd__inv_2 _14110_ (.A(_07030_),
    .Y(_00305_));
 sky130_fd_sc_hd__inv_2 _14111_ (.A(_07030_),
    .Y(_00306_));
 sky130_fd_sc_hd__inv_2 _14112_ (.A(_07030_),
    .Y(_00307_));
 sky130_fd_sc_hd__inv_2 _14113_ (.A(_07030_),
    .Y(_00308_));
 sky130_fd_sc_hd__clkbuf_8 _14114_ (.A(_04755_),
    .X(_07031_));
 sky130_fd_sc_hd__inv_2 _14115_ (.A(_07031_),
    .Y(_00309_));
 sky130_fd_sc_hd__inv_2 _14116_ (.A(_07031_),
    .Y(_00310_));
 sky130_fd_sc_hd__inv_2 _14117_ (.A(_07031_),
    .Y(_00311_));
 sky130_fd_sc_hd__inv_2 _14118_ (.A(_07031_),
    .Y(_00312_));
 sky130_fd_sc_hd__inv_2 _14119_ (.A(_07031_),
    .Y(_00313_));
 sky130_fd_sc_hd__inv_2 _14120_ (.A(_07031_),
    .Y(_00314_));
 sky130_fd_sc_hd__inv_2 _14121_ (.A(_07031_),
    .Y(_00315_));
 sky130_fd_sc_hd__inv_2 _14122_ (.A(_07031_),
    .Y(_00316_));
 sky130_fd_sc_hd__inv_2 _14123_ (.A(_07031_),
    .Y(_00317_));
 sky130_fd_sc_hd__inv_2 _14124_ (.A(_07031_),
    .Y(_00318_));
 sky130_fd_sc_hd__dfxtp_1 _14125_ (.CLK(clknet_leaf_106_clk),
    .D(_00319_),
    .Q(\regs[9][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14126_ (.CLK(clknet_leaf_131_clk),
    .D(_00320_),
    .Q(\regs[9][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14127_ (.CLK(clknet_leaf_129_clk),
    .D(_00321_),
    .Q(\regs[9][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14128_ (.CLK(clknet_leaf_135_clk),
    .D(_00322_),
    .Q(\regs[9][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14129_ (.CLK(clknet_leaf_128_clk),
    .D(_00323_),
    .Q(\regs[9][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14130_ (.CLK(clknet_leaf_133_clk),
    .D(_00324_),
    .Q(\regs[9][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14131_ (.CLK(clknet_leaf_105_clk),
    .D(_00325_),
    .Q(\regs[9][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14132_ (.CLK(clknet_leaf_126_clk),
    .D(_00326_),
    .Q(\regs[9][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14133_ (.CLK(clknet_leaf_133_clk),
    .D(_00327_),
    .Q(\regs[9][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14134_ (.CLK(clknet_leaf_104_clk),
    .D(_00328_),
    .Q(\regs[9][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14135_ (.CLK(clknet_leaf_104_clk),
    .D(_00329_),
    .Q(\regs[9][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14136_ (.CLK(clknet_leaf_98_clk),
    .D(_00330_),
    .Q(\regs[9][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14137_ (.CLK(clknet_leaf_97_clk),
    .D(_00331_),
    .Q(\regs[9][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14138_ (.CLK(clknet_leaf_101_clk),
    .D(_00332_),
    .Q(\regs[9][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14139_ (.CLK(clknet_leaf_97_clk),
    .D(_00333_),
    .Q(\regs[9][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14140_ (.CLK(clknet_leaf_104_clk),
    .D(_00334_),
    .Q(\regs[9][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14141_ (.CLK(clknet_leaf_98_clk),
    .D(_00335_),
    .Q(\regs[9][16] ));
 sky130_fd_sc_hd__dfxtp_1 _14142_ (.CLK(clknet_leaf_103_clk),
    .D(_00336_),
    .Q(\regs[9][17] ));
 sky130_fd_sc_hd__dfxtp_1 _14143_ (.CLK(clknet_leaf_101_clk),
    .D(_00337_),
    .Q(\regs[9][18] ));
 sky130_fd_sc_hd__dfxtp_1 _14144_ (.CLK(clknet_leaf_102_clk),
    .D(_00338_),
    .Q(\regs[9][19] ));
 sky130_fd_sc_hd__dfxtp_1 _14145_ (.CLK(clknet_leaf_7_clk),
    .D(_00339_),
    .Q(\regs[9][20] ));
 sky130_fd_sc_hd__dfxtp_1 _14146_ (.CLK(clknet_leaf_65_clk),
    .D(_00340_),
    .Q(\regs[9][21] ));
 sky130_fd_sc_hd__dfxtp_1 _14147_ (.CLK(clknet_leaf_66_clk),
    .D(_00341_),
    .Q(\regs[9][22] ));
 sky130_fd_sc_hd__dfxtp_1 _14148_ (.CLK(clknet_leaf_27_clk),
    .D(_00342_),
    .Q(\regs[9][23] ));
 sky130_fd_sc_hd__dfxtp_1 _14149_ (.CLK(clknet_leaf_20_clk),
    .D(_00343_),
    .Q(\regs[9][24] ));
 sky130_fd_sc_hd__dfxtp_1 _14150_ (.CLK(clknet_leaf_7_clk),
    .D(_00344_),
    .Q(\regs[9][25] ));
 sky130_fd_sc_hd__dfxtp_1 _14151_ (.CLK(clknet_leaf_66_clk),
    .D(_00345_),
    .Q(\regs[9][26] ));
 sky130_fd_sc_hd__dfxtp_1 _14152_ (.CLK(clknet_leaf_65_clk),
    .D(_00346_),
    .Q(\regs[9][27] ));
 sky130_fd_sc_hd__dfxtp_1 _14153_ (.CLK(clknet_leaf_7_clk),
    .D(_00347_),
    .Q(\regs[9][28] ));
 sky130_fd_sc_hd__dfxtp_1 _14154_ (.CLK(clknet_leaf_21_clk),
    .D(_00348_),
    .Q(\regs[9][29] ));
 sky130_fd_sc_hd__dfxtp_1 _14155_ (.CLK(clknet_leaf_115_clk),
    .D(_00349_),
    .Q(\regs[9][30] ));
 sky130_fd_sc_hd__dfxtp_1 _14156_ (.CLK(clknet_leaf_112_clk),
    .D(_00350_),
    .Q(\regs[9][31] ));
 sky130_fd_sc_hd__dfxtp_1 _14157_ (.CLK(clknet_leaf_125_clk),
    .D(_00351_),
    .Q(\regs[7][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14158_ (.CLK(clknet_leaf_134_clk),
    .D(_00352_),
    .Q(\regs[7][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14159_ (.CLK(clknet_leaf_129_clk),
    .D(_00353_),
    .Q(\regs[7][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14160_ (.CLK(clknet_leaf_0_clk),
    .D(_00354_),
    .Q(\regs[7][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14161_ (.CLK(clknet_leaf_130_clk),
    .D(_00355_),
    .Q(\regs[7][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14162_ (.CLK(clknet_leaf_0_clk),
    .D(_00356_),
    .Q(\regs[7][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14163_ (.CLK(clknet_leaf_105_clk),
    .D(_00357_),
    .Q(\regs[7][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14164_ (.CLK(clknet_leaf_127_clk),
    .D(_00358_),
    .Q(\regs[7][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14165_ (.CLK(clknet_leaf_1_clk),
    .D(_00359_),
    .Q(\regs[7][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14166_ (.CLK(clknet_leaf_125_clk),
    .D(_00360_),
    .Q(\regs[7][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14167_ (.CLK(clknet_leaf_110_clk),
    .D(_00361_),
    .Q(\regs[7][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14168_ (.CLK(clknet_leaf_96_clk),
    .D(_00362_),
    .Q(\regs[7][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14169_ (.CLK(clknet_leaf_98_clk),
    .D(_00363_),
    .Q(\regs[7][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14170_ (.CLK(clknet_leaf_90_clk),
    .D(_00364_),
    .Q(\regs[7][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14171_ (.CLK(clknet_leaf_95_clk),
    .D(_00365_),
    .Q(\regs[7][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14172_ (.CLK(clknet_leaf_109_clk),
    .D(_00366_),
    .Q(\regs[7][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14173_ (.CLK(clknet_leaf_91_clk),
    .D(_00367_),
    .Q(\regs[7][16] ));
 sky130_fd_sc_hd__dfxtp_1 _14174_ (.CLK(clknet_leaf_100_clk),
    .D(_00368_),
    .Q(\regs[7][17] ));
 sky130_fd_sc_hd__dfxtp_1 _14175_ (.CLK(clknet_leaf_111_clk),
    .D(_00369_),
    .Q(\regs[7][18] ));
 sky130_fd_sc_hd__dfxtp_1 _14176_ (.CLK(clknet_leaf_91_clk),
    .D(_00370_),
    .Q(\regs[7][19] ));
 sky130_fd_sc_hd__dfxtp_1 _14177_ (.CLK(clknet_leaf_8_clk),
    .D(_00371_),
    .Q(\regs[7][20] ));
 sky130_fd_sc_hd__dfxtp_1 _14178_ (.CLK(clknet_leaf_63_clk),
    .D(_00372_),
    .Q(\regs[7][21] ));
 sky130_fd_sc_hd__dfxtp_1 _14179_ (.CLK(clknet_leaf_64_clk),
    .D(_00373_),
    .Q(\regs[7][22] ));
 sky130_fd_sc_hd__dfxtp_1 _14180_ (.CLK(clknet_leaf_28_clk),
    .D(_00374_),
    .Q(\regs[7][23] ));
 sky130_fd_sc_hd__dfxtp_1 _14181_ (.CLK(clknet_leaf_25_clk),
    .D(_00375_),
    .Q(\regs[7][24] ));
 sky130_fd_sc_hd__dfxtp_1 _14182_ (.CLK(clknet_leaf_9_clk),
    .D(_00376_),
    .Q(\regs[7][25] ));
 sky130_fd_sc_hd__dfxtp_1 _14183_ (.CLK(clknet_leaf_69_clk),
    .D(_00377_),
    .Q(\regs[7][26] ));
 sky130_fd_sc_hd__dfxtp_1 _14184_ (.CLK(clknet_leaf_66_clk),
    .D(_00378_),
    .Q(\regs[7][27] ));
 sky130_fd_sc_hd__dfxtp_1 _14185_ (.CLK(clknet_leaf_8_clk),
    .D(_00379_),
    .Q(\regs[7][28] ));
 sky130_fd_sc_hd__dfxtp_1 _14186_ (.CLK(clknet_leaf_56_clk),
    .D(_00380_),
    .Q(\regs[7][29] ));
 sky130_fd_sc_hd__dfxtp_1 _14187_ (.CLK(clknet_leaf_116_clk),
    .D(_00381_),
    .Q(\regs[7][30] ));
 sky130_fd_sc_hd__dfxtp_1 _14188_ (.CLK(clknet_leaf_74_clk),
    .D(_00382_),
    .Q(\regs[7][31] ));
 sky130_fd_sc_hd__dfxtp_1 _14189_ (.CLK(clknet_leaf_126_clk),
    .D(_00383_),
    .Q(\regs[10][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14190_ (.CLK(clknet_leaf_132_clk),
    .D(_00384_),
    .Q(\regs[10][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14191_ (.CLK(clknet_leaf_128_clk),
    .D(_00385_),
    .Q(\regs[10][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14192_ (.CLK(clknet_leaf_135_clk),
    .D(_00386_),
    .Q(\regs[10][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14193_ (.CLK(clknet_leaf_128_clk),
    .D(_00387_),
    .Q(\regs[10][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14194_ (.CLK(clknet_leaf_133_clk),
    .D(_00388_),
    .Q(\regs[10][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14195_ (.CLK(clknet_leaf_105_clk),
    .D(_00389_),
    .Q(\regs[10][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14196_ (.CLK(clknet_leaf_126_clk),
    .D(_00390_),
    .Q(\regs[10][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14197_ (.CLK(clknet_leaf_135_clk),
    .D(_00391_),
    .Q(\regs[10][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14198_ (.CLK(clknet_leaf_105_clk),
    .D(_00392_),
    .Q(\regs[10][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14199_ (.CLK(clknet_leaf_103_clk),
    .D(_00393_),
    .Q(\regs[10][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14200_ (.CLK(clknet_leaf_98_clk),
    .D(_00394_),
    .Q(\regs[10][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14201_ (.CLK(clknet_leaf_102_clk),
    .D(_00395_),
    .Q(\regs[10][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14202_ (.CLK(clknet_leaf_101_clk),
    .D(_00396_),
    .Q(\regs[10][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14203_ (.CLK(clknet_leaf_97_clk),
    .D(_00397_),
    .Q(\regs[10][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14204_ (.CLK(clknet_leaf_106_clk),
    .D(_00398_),
    .Q(\regs[10][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14205_ (.CLK(clknet_leaf_97_clk),
    .D(_00399_),
    .Q(\regs[10][16] ));
 sky130_fd_sc_hd__dfxtp_1 _14206_ (.CLK(clknet_leaf_103_clk),
    .D(_00400_),
    .Q(\regs[10][17] ));
 sky130_fd_sc_hd__dfxtp_1 _14207_ (.CLK(clknet_leaf_101_clk),
    .D(_00401_),
    .Q(\regs[10][18] ));
 sky130_fd_sc_hd__dfxtp_1 _14208_ (.CLK(clknet_leaf_103_clk),
    .D(_00402_),
    .Q(\regs[10][19] ));
 sky130_fd_sc_hd__dfxtp_1 _14209_ (.CLK(clknet_leaf_6_clk),
    .D(_00403_),
    .Q(\regs[10][20] ));
 sky130_fd_sc_hd__dfxtp_1 _14210_ (.CLK(clknet_leaf_65_clk),
    .D(_00404_),
    .Q(\regs[10][21] ));
 sky130_fd_sc_hd__dfxtp_1 _14211_ (.CLK(clknet_leaf_65_clk),
    .D(_00405_),
    .Q(\regs[10][22] ));
 sky130_fd_sc_hd__dfxtp_1 _14212_ (.CLK(clknet_leaf_28_clk),
    .D(_00406_),
    .Q(\regs[10][23] ));
 sky130_fd_sc_hd__dfxtp_1 _14213_ (.CLK(clknet_leaf_20_clk),
    .D(_00407_),
    .Q(\regs[10][24] ));
 sky130_fd_sc_hd__dfxtp_1 _14214_ (.CLK(clknet_leaf_6_clk),
    .D(_00408_),
    .Q(\regs[10][25] ));
 sky130_fd_sc_hd__dfxtp_1 _14215_ (.CLK(clknet_leaf_69_clk),
    .D(_00409_),
    .Q(\regs[10][26] ));
 sky130_fd_sc_hd__dfxtp_1 _14216_ (.CLK(clknet_leaf_65_clk),
    .D(_00410_),
    .Q(\regs[10][27] ));
 sky130_fd_sc_hd__dfxtp_1 _14217_ (.CLK(clknet_leaf_7_clk),
    .D(_00411_),
    .Q(\regs[10][28] ));
 sky130_fd_sc_hd__dfxtp_1 _14218_ (.CLK(clknet_leaf_21_clk),
    .D(_00412_),
    .Q(\regs[10][29] ));
 sky130_fd_sc_hd__dfxtp_1 _14219_ (.CLK(clknet_leaf_114_clk),
    .D(_00413_),
    .Q(\regs[10][30] ));
 sky130_fd_sc_hd__dfxtp_1 _14220_ (.CLK(clknet_leaf_115_clk),
    .D(_00414_),
    .Q(\regs[10][31] ));
 sky130_fd_sc_hd__dfxtp_1 _14221_ (.CLK(clknet_leaf_125_clk),
    .D(_00415_),
    .Q(\regs[12][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14222_ (.CLK(clknet_leaf_134_clk),
    .D(_00416_),
    .Q(\regs[12][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14223_ (.CLK(clknet_leaf_129_clk),
    .D(_00417_),
    .Q(\regs[12][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14224_ (.CLK(clknet_leaf_133_clk),
    .D(_00418_),
    .Q(\regs[12][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14225_ (.CLK(clknet_leaf_128_clk),
    .D(_00419_),
    .Q(\regs[12][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14226_ (.CLK(clknet_leaf_3_clk),
    .D(_00420_),
    .Q(\regs[12][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14227_ (.CLK(clknet_leaf_106_clk),
    .D(_00421_),
    .Q(\regs[12][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14228_ (.CLK(clknet_leaf_126_clk),
    .D(_00422_),
    .Q(\regs[12][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14229_ (.CLK(clknet_leaf_133_clk),
    .D(_00423_),
    .Q(\regs[12][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14230_ (.CLK(clknet_leaf_104_clk),
    .D(_00424_),
    .Q(\regs[12][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14231_ (.CLK(clknet_leaf_104_clk),
    .D(_00425_),
    .Q(\regs[12][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14232_ (.CLK(clknet_leaf_96_clk),
    .D(_00426_),
    .Q(\regs[12][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14233_ (.CLK(clknet_leaf_102_clk),
    .D(_00427_),
    .Q(\regs[12][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14234_ (.CLK(clknet_leaf_90_clk),
    .D(_00428_),
    .Q(\regs[12][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14235_ (.CLK(clknet_leaf_99_clk),
    .D(_00429_),
    .Q(\regs[12][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14236_ (.CLK(clknet_leaf_110_clk),
    .D(_00430_),
    .Q(\regs[12][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14237_ (.CLK(clknet_leaf_91_clk),
    .D(_00431_),
    .Q(\regs[12][16] ));
 sky130_fd_sc_hd__dfxtp_1 _14238_ (.CLK(clknet_leaf_99_clk),
    .D(_00432_),
    .Q(\regs[12][17] ));
 sky130_fd_sc_hd__dfxtp_1 _14239_ (.CLK(clknet_leaf_100_clk),
    .D(_00433_),
    .Q(\regs[12][18] ));
 sky130_fd_sc_hd__dfxtp_1 _14240_ (.CLK(clknet_leaf_91_clk),
    .D(_00434_),
    .Q(\regs[12][19] ));
 sky130_fd_sc_hd__dfxtp_1 _14241_ (.CLK(clknet_leaf_10_clk),
    .D(_00435_),
    .Q(\regs[12][20] ));
 sky130_fd_sc_hd__dfxtp_1 _14242_ (.CLK(clknet_leaf_81_clk),
    .D(_00436_),
    .Q(\regs[12][21] ));
 sky130_fd_sc_hd__dfxtp_1 _14243_ (.CLK(clknet_leaf_64_clk),
    .D(_00437_),
    .Q(\regs[12][22] ));
 sky130_fd_sc_hd__dfxtp_1 _14244_ (.CLK(clknet_leaf_25_clk),
    .D(_00438_),
    .Q(\regs[12][23] ));
 sky130_fd_sc_hd__dfxtp_1 _14245_ (.CLK(clknet_leaf_19_clk),
    .D(_00439_),
    .Q(\regs[12][24] ));
 sky130_fd_sc_hd__dfxtp_1 _14246_ (.CLK(clknet_leaf_10_clk),
    .D(_00440_),
    .Q(\regs[12][25] ));
 sky130_fd_sc_hd__dfxtp_1 _14247_ (.CLK(clknet_leaf_70_clk),
    .D(_00441_),
    .Q(\regs[12][26] ));
 sky130_fd_sc_hd__dfxtp_1 _14248_ (.CLK(clknet_leaf_64_clk),
    .D(_00442_),
    .Q(\regs[12][27] ));
 sky130_fd_sc_hd__dfxtp_1 _14249_ (.CLK(clknet_leaf_10_clk),
    .D(_00443_),
    .Q(\regs[12][28] ));
 sky130_fd_sc_hd__dfxtp_1 _14250_ (.CLK(clknet_leaf_71_clk),
    .D(_00444_),
    .Q(\regs[12][29] ));
 sky130_fd_sc_hd__dfxtp_1 _14251_ (.CLK(clknet_leaf_112_clk),
    .D(_00445_),
    .Q(\regs[12][30] ));
 sky130_fd_sc_hd__dfxtp_1 _14252_ (.CLK(clknet_leaf_74_clk),
    .D(_00446_),
    .Q(\regs[12][31] ));
 sky130_fd_sc_hd__dfxtp_1 _14253_ (.CLK(clknet_leaf_128_clk),
    .D(_00447_),
    .Q(\regs[15][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14254_ (.CLK(clknet_leaf_133_clk),
    .D(_00448_),
    .Q(\regs[15][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14255_ (.CLK(clknet_leaf_130_clk),
    .D(_00449_),
    .Q(\regs[15][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14256_ (.CLK(clknet_leaf_133_clk),
    .D(_00450_),
    .Q(\regs[15][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14257_ (.CLK(clknet_leaf_130_clk),
    .D(_00451_),
    .Q(\regs[15][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14258_ (.CLK(clknet_leaf_2_clk),
    .D(_00452_),
    .Q(\regs[15][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14259_ (.CLK(clknet_leaf_106_clk),
    .D(_00453_),
    .Q(\regs[15][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14260_ (.CLK(clknet_leaf_127_clk),
    .D(_00454_),
    .Q(\regs[15][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14261_ (.CLK(clknet_leaf_2_clk),
    .D(_00455_),
    .Q(\regs[15][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14262_ (.CLK(clknet_leaf_106_clk),
    .D(_00456_),
    .Q(\regs[15][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14263_ (.CLK(clknet_leaf_104_clk),
    .D(_00457_),
    .Q(\regs[15][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14264_ (.CLK(clknet_leaf_96_clk),
    .D(_00458_),
    .Q(\regs[15][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14265_ (.CLK(clknet_leaf_104_clk),
    .D(_00459_),
    .Q(\regs[15][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14266_ (.CLK(clknet_leaf_90_clk),
    .D(_00460_),
    .Q(\regs[15][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14267_ (.CLK(clknet_leaf_98_clk),
    .D(_00461_),
    .Q(\regs[15][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14268_ (.CLK(clknet_leaf_107_clk),
    .D(_00462_),
    .Q(\regs[15][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14269_ (.CLK(clknet_leaf_99_clk),
    .D(_00463_),
    .Q(\regs[15][16] ));
 sky130_fd_sc_hd__dfxtp_1 _14270_ (.CLK(clknet_leaf_99_clk),
    .D(_00464_),
    .Q(\regs[15][17] ));
 sky130_fd_sc_hd__dfxtp_1 _14271_ (.CLK(clknet_leaf_100_clk),
    .D(_00465_),
    .Q(\regs[15][18] ));
 sky130_fd_sc_hd__dfxtp_1 _14272_ (.CLK(clknet_leaf_90_clk),
    .D(_00466_),
    .Q(\regs[15][19] ));
 sky130_fd_sc_hd__dfxtp_1 _14273_ (.CLK(clknet_leaf_9_clk),
    .D(_00467_),
    .Q(\regs[15][20] ));
 sky130_fd_sc_hd__dfxtp_1 _14274_ (.CLK(clknet_leaf_81_clk),
    .D(_00468_),
    .Q(\regs[15][21] ));
 sky130_fd_sc_hd__dfxtp_1 _14275_ (.CLK(clknet_leaf_65_clk),
    .D(_00469_),
    .Q(\regs[15][22] ));
 sky130_fd_sc_hd__dfxtp_1 _14276_ (.CLK(clknet_leaf_27_clk),
    .D(_00470_),
    .Q(\regs[15][23] ));
 sky130_fd_sc_hd__dfxtp_1 _14277_ (.CLK(clknet_leaf_19_clk),
    .D(_00471_),
    .Q(\regs[15][24] ));
 sky130_fd_sc_hd__dfxtp_1 _14278_ (.CLK(clknet_leaf_9_clk),
    .D(_00472_),
    .Q(\regs[15][25] ));
 sky130_fd_sc_hd__dfxtp_1 _14279_ (.CLK(clknet_leaf_69_clk),
    .D(_00473_),
    .Q(\regs[15][26] ));
 sky130_fd_sc_hd__dfxtp_1 _14280_ (.CLK(clknet_leaf_65_clk),
    .D(_00474_),
    .Q(\regs[15][27] ));
 sky130_fd_sc_hd__dfxtp_1 _14281_ (.CLK(clknet_leaf_9_clk),
    .D(_00475_),
    .Q(\regs[15][28] ));
 sky130_fd_sc_hd__dfxtp_1 _14282_ (.CLK(clknet_leaf_70_clk),
    .D(_00476_),
    .Q(\regs[15][29] ));
 sky130_fd_sc_hd__dfxtp_1 _14283_ (.CLK(clknet_leaf_115_clk),
    .D(_00477_),
    .Q(\regs[15][30] ));
 sky130_fd_sc_hd__dfxtp_1 _14284_ (.CLK(clknet_leaf_74_clk),
    .D(_00478_),
    .Q(\regs[15][31] ));
 sky130_fd_sc_hd__dfxtp_1 _14285_ (.CLK(clknet_leaf_125_clk),
    .D(_00479_),
    .Q(\regs[5][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14286_ (.CLK(clknet_leaf_130_clk),
    .D(_00480_),
    .Q(\regs[5][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14287_ (.CLK(clknet_leaf_129_clk),
    .D(_00481_),
    .Q(\regs[5][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14288_ (.CLK(clknet_leaf_135_clk),
    .D(_00482_),
    .Q(\regs[5][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14289_ (.CLK(clknet_leaf_131_clk),
    .D(_00483_),
    .Q(\regs[5][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14290_ (.CLK(clknet_leaf_1_clk),
    .D(_00484_),
    .Q(\regs[5][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14291_ (.CLK(clknet_leaf_105_clk),
    .D(_00485_),
    .Q(\regs[5][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14292_ (.CLK(clknet_leaf_127_clk),
    .D(_00486_),
    .Q(\regs[5][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14293_ (.CLK(clknet_leaf_1_clk),
    .D(_00487_),
    .Q(\regs[5][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14294_ (.CLK(clknet_leaf_106_clk),
    .D(_00488_),
    .Q(\regs[5][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14295_ (.CLK(clknet_leaf_110_clk),
    .D(_00489_),
    .Q(\regs[5][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14296_ (.CLK(clknet_leaf_95_clk),
    .D(_00490_),
    .Q(\regs[5][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14297_ (.CLK(clknet_leaf_97_clk),
    .D(_00491_),
    .Q(\regs[5][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14298_ (.CLK(clknet_leaf_92_clk),
    .D(_00492_),
    .Q(\regs[5][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14299_ (.CLK(clknet_leaf_94_clk),
    .D(_00493_),
    .Q(\regs[5][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14300_ (.CLK(clknet_leaf_110_clk),
    .D(_00494_),
    .Q(\regs[5][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14301_ (.CLK(clknet_leaf_94_clk),
    .D(_00495_),
    .Q(\regs[5][16] ));
 sky130_fd_sc_hd__dfxtp_1 _14302_ (.CLK(clknet_leaf_100_clk),
    .D(_00496_),
    .Q(\regs[5][17] ));
 sky130_fd_sc_hd__dfxtp_1 _14303_ (.CLK(clknet_leaf_100_clk),
    .D(_00497_),
    .Q(\regs[5][18] ));
 sky130_fd_sc_hd__dfxtp_1 _14304_ (.CLK(clknet_leaf_91_clk),
    .D(_00498_),
    .Q(\regs[5][19] ));
 sky130_fd_sc_hd__dfxtp_1 _14305_ (.CLK(clknet_leaf_8_clk),
    .D(_00499_),
    .Q(\regs[5][20] ));
 sky130_fd_sc_hd__dfxtp_1 _14306_ (.CLK(clknet_leaf_63_clk),
    .D(_00500_),
    .Q(\regs[5][21] ));
 sky130_fd_sc_hd__dfxtp_1 _14307_ (.CLK(clknet_leaf_62_clk),
    .D(_00501_),
    .Q(\regs[5][22] ));
 sky130_fd_sc_hd__dfxtp_1 _14308_ (.CLK(clknet_leaf_29_clk),
    .D(_00502_),
    .Q(\regs[5][23] ));
 sky130_fd_sc_hd__dfxtp_1 _14309_ (.CLK(clknet_leaf_22_clk),
    .D(_00503_),
    .Q(\regs[5][24] ));
 sky130_fd_sc_hd__dfxtp_1 _14310_ (.CLK(clknet_leaf_9_clk),
    .D(_00504_),
    .Q(\regs[5][25] ));
 sky130_fd_sc_hd__dfxtp_1 _14311_ (.CLK(clknet_leaf_69_clk),
    .D(_00505_),
    .Q(\regs[5][26] ));
 sky130_fd_sc_hd__dfxtp_1 _14312_ (.CLK(clknet_leaf_64_clk),
    .D(_00506_),
    .Q(\regs[5][27] ));
 sky130_fd_sc_hd__dfxtp_1 _14313_ (.CLK(clknet_leaf_8_clk),
    .D(_00507_),
    .Q(\regs[5][28] ));
 sky130_fd_sc_hd__dfxtp_1 _14314_ (.CLK(clknet_leaf_71_clk),
    .D(_00508_),
    .Q(\regs[5][29] ));
 sky130_fd_sc_hd__dfxtp_1 _14315_ (.CLK(clknet_leaf_73_clk),
    .D(_00509_),
    .Q(\regs[5][30] ));
 sky130_fd_sc_hd__dfxtp_1 _14316_ (.CLK(clknet_leaf_74_clk),
    .D(_00510_),
    .Q(\regs[5][31] ));
 sky130_fd_sc_hd__dfxtp_1 _14317_ (.CLK(clknet_leaf_126_clk),
    .D(_00511_),
    .Q(\regs[8][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14318_ (.CLK(clknet_leaf_134_clk),
    .D(_00512_),
    .Q(\regs[8][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14319_ (.CLK(clknet_leaf_128_clk),
    .D(_00513_),
    .Q(\regs[8][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14320_ (.CLK(clknet_leaf_133_clk),
    .D(_00514_),
    .Q(\regs[8][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14321_ (.CLK(clknet_leaf_127_clk),
    .D(_00515_),
    .Q(\regs[8][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14322_ (.CLK(clknet_leaf_133_clk),
    .D(_00516_),
    .Q(\regs[8][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14323_ (.CLK(clknet_leaf_105_clk),
    .D(_00517_),
    .Q(\regs[8][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14324_ (.CLK(clknet_leaf_126_clk),
    .D(_00518_),
    .Q(\regs[8][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14325_ (.CLK(clknet_leaf_133_clk),
    .D(_00519_),
    .Q(\regs[8][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14326_ (.CLK(clknet_leaf_104_clk),
    .D(_00520_),
    .Q(\regs[8][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14327_ (.CLK(clknet_leaf_104_clk),
    .D(_00521_),
    .Q(\regs[8][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14328_ (.CLK(clknet_leaf_98_clk),
    .D(_00522_),
    .Q(\regs[8][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14329_ (.CLK(clknet_leaf_97_clk),
    .D(_00523_),
    .Q(\regs[8][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14330_ (.CLK(clknet_leaf_102_clk),
    .D(_00524_),
    .Q(\regs[8][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14331_ (.CLK(clknet_leaf_96_clk),
    .D(_00525_),
    .Q(\regs[8][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14332_ (.CLK(clknet_leaf_104_clk),
    .D(_00526_),
    .Q(\regs[8][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14333_ (.CLK(clknet_leaf_96_clk),
    .D(_00527_),
    .Q(\regs[8][16] ));
 sky130_fd_sc_hd__dfxtp_1 _14334_ (.CLK(clknet_leaf_103_clk),
    .D(_00528_),
    .Q(\regs[8][17] ));
 sky130_fd_sc_hd__dfxtp_1 _14335_ (.CLK(clknet_leaf_101_clk),
    .D(_00529_),
    .Q(\regs[8][18] ));
 sky130_fd_sc_hd__dfxtp_1 _14336_ (.CLK(clknet_leaf_102_clk),
    .D(_00530_),
    .Q(\regs[8][19] ));
 sky130_fd_sc_hd__dfxtp_1 _14337_ (.CLK(clknet_leaf_6_clk),
    .D(_00531_),
    .Q(\regs[8][20] ));
 sky130_fd_sc_hd__dfxtp_1 _14338_ (.CLK(clknet_leaf_81_clk),
    .D(_00532_),
    .Q(\regs[8][21] ));
 sky130_fd_sc_hd__dfxtp_1 _14339_ (.CLK(clknet_leaf_66_clk),
    .D(_00533_),
    .Q(\regs[8][22] ));
 sky130_fd_sc_hd__dfxtp_1 _14340_ (.CLK(clknet_leaf_25_clk),
    .D(_00534_),
    .Q(\regs[8][23] ));
 sky130_fd_sc_hd__dfxtp_1 _14341_ (.CLK(clknet_leaf_20_clk),
    .D(_00535_),
    .Q(\regs[8][24] ));
 sky130_fd_sc_hd__dfxtp_1 _14342_ (.CLK(clknet_leaf_12_clk),
    .D(_00536_),
    .Q(\regs[8][25] ));
 sky130_fd_sc_hd__dfxtp_1 _14343_ (.CLK(clknet_leaf_66_clk),
    .D(_00537_),
    .Q(\regs[8][26] ));
 sky130_fd_sc_hd__dfxtp_1 _14344_ (.CLK(clknet_leaf_65_clk),
    .D(_00538_),
    .Q(\regs[8][27] ));
 sky130_fd_sc_hd__dfxtp_1 _14345_ (.CLK(clknet_leaf_7_clk),
    .D(_00539_),
    .Q(\regs[8][28] ));
 sky130_fd_sc_hd__dfxtp_1 _14346_ (.CLK(clknet_leaf_20_clk),
    .D(_00540_),
    .Q(\regs[8][29] ));
 sky130_fd_sc_hd__dfxtp_1 _14347_ (.CLK(clknet_leaf_115_clk),
    .D(_00541_),
    .Q(\regs[8][30] ));
 sky130_fd_sc_hd__dfxtp_1 _14348_ (.CLK(clknet_leaf_77_clk),
    .D(_00542_),
    .Q(\regs[8][31] ));
 sky130_fd_sc_hd__dfstp_1 _14349_ (.CLK(clknet_leaf_56_clk),
    .D(_00000_),
    .SET_B(_00068_),
    .Q(\core_state[0] ));
 sky130_fd_sc_hd__dfrtp_4 _14350_ (.CLK(clknet_leaf_57_clk),
    .D(_00001_),
    .RESET_B(_00069_),
    .Q(\core_state[1] ));
 sky130_fd_sc_hd__dfrtp_1 _14351_ (.CLK(clknet_leaf_56_clk),
    .D(_00002_),
    .RESET_B(_00070_),
    .Q(\core_state[2] ));
 sky130_fd_sc_hd__dfrtp_1 _14352_ (.CLK(clknet_leaf_56_clk),
    .D(_00003_),
    .RESET_B(_00071_),
    .Q(\core_state[3] ));
 sky130_fd_sc_hd__dfxtp_1 _14353_ (.CLK(clknet_leaf_127_clk),
    .D(_00543_),
    .Q(\regs[13][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14354_ (.CLK(clknet_leaf_133_clk),
    .D(_00544_),
    .Q(\regs[13][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14355_ (.CLK(clknet_leaf_130_clk),
    .D(_00545_),
    .Q(\regs[13][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14356_ (.CLK(clknet_leaf_133_clk),
    .D(_00546_),
    .Q(\regs[13][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14357_ (.CLK(clknet_leaf_128_clk),
    .D(_00547_),
    .Q(\regs[13][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14358_ (.CLK(clknet_leaf_2_clk),
    .D(_00548_),
    .Q(\regs[13][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14359_ (.CLK(clknet_leaf_105_clk),
    .D(_00549_),
    .Q(\regs[13][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14360_ (.CLK(clknet_leaf_126_clk),
    .D(_00550_),
    .Q(\regs[13][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14361_ (.CLK(clknet_leaf_132_clk),
    .D(_00551_),
    .Q(\regs[13][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14362_ (.CLK(clknet_leaf_106_clk),
    .D(_00552_),
    .Q(\regs[13][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14363_ (.CLK(clknet_leaf_101_clk),
    .D(_00553_),
    .Q(\regs[13][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14364_ (.CLK(clknet_leaf_96_clk),
    .D(_00554_),
    .Q(\regs[13][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14365_ (.CLK(clknet_leaf_102_clk),
    .D(_00555_),
    .Q(\regs[13][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14366_ (.CLK(clknet_leaf_91_clk),
    .D(_00556_),
    .Q(\regs[13][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14367_ (.CLK(clknet_leaf_98_clk),
    .D(_00557_),
    .Q(\regs[13][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14368_ (.CLK(clknet_leaf_101_clk),
    .D(_00558_),
    .Q(\regs[13][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14369_ (.CLK(clknet_leaf_91_clk),
    .D(_00559_),
    .Q(\regs[13][16] ));
 sky130_fd_sc_hd__dfxtp_1 _14370_ (.CLK(clknet_leaf_99_clk),
    .D(_00560_),
    .Q(\regs[13][17] ));
 sky130_fd_sc_hd__dfxtp_1 _14371_ (.CLK(clknet_leaf_100_clk),
    .D(_00561_),
    .Q(\regs[13][18] ));
 sky130_fd_sc_hd__dfxtp_1 _14372_ (.CLK(clknet_leaf_91_clk),
    .D(_00562_),
    .Q(\regs[13][19] ));
 sky130_fd_sc_hd__dfxtp_1 _14373_ (.CLK(clknet_leaf_9_clk),
    .D(_00563_),
    .Q(\regs[13][20] ));
 sky130_fd_sc_hd__dfxtp_1 _14374_ (.CLK(clknet_leaf_81_clk),
    .D(_00564_),
    .Q(\regs[13][21] ));
 sky130_fd_sc_hd__dfxtp_1 _14375_ (.CLK(clknet_leaf_64_clk),
    .D(_00565_),
    .Q(\regs[13][22] ));
 sky130_fd_sc_hd__dfxtp_1 _14376_ (.CLK(clknet_leaf_27_clk),
    .D(_00566_),
    .Q(\regs[13][23] ));
 sky130_fd_sc_hd__dfxtp_1 _14377_ (.CLK(clknet_leaf_19_clk),
    .D(_00567_),
    .Q(\regs[13][24] ));
 sky130_fd_sc_hd__dfxtp_1 _14378_ (.CLK(clknet_leaf_10_clk),
    .D(_00568_),
    .Q(\regs[13][25] ));
 sky130_fd_sc_hd__dfxtp_1 _14379_ (.CLK(clknet_leaf_70_clk),
    .D(_00569_),
    .Q(\regs[13][26] ));
 sky130_fd_sc_hd__dfxtp_1 _14380_ (.CLK(clknet_leaf_64_clk),
    .D(_00570_),
    .Q(\regs[13][27] ));
 sky130_fd_sc_hd__dfxtp_1 _14381_ (.CLK(clknet_leaf_10_clk),
    .D(_00571_),
    .Q(\regs[13][28] ));
 sky130_fd_sc_hd__dfxtp_1 _14382_ (.CLK(clknet_leaf_70_clk),
    .D(_00572_),
    .Q(\regs[13][29] ));
 sky130_fd_sc_hd__dfxtp_1 _14383_ (.CLK(clknet_leaf_112_clk),
    .D(_00573_),
    .Q(\regs[13][30] ));
 sky130_fd_sc_hd__dfxtp_1 _14384_ (.CLK(clknet_leaf_74_clk),
    .D(_00574_),
    .Q(\regs[13][31] ));
 sky130_fd_sc_hd__dfxtp_1 _14385_ (.CLK(clknet_leaf_127_clk),
    .D(_00575_),
    .Q(\regs[14][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14386_ (.CLK(clknet_leaf_134_clk),
    .D(_00576_),
    .Q(\regs[14][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14387_ (.CLK(clknet_leaf_130_clk),
    .D(_00577_),
    .Q(\regs[14][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14388_ (.CLK(clknet_leaf_133_clk),
    .D(_00578_),
    .Q(\regs[14][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14389_ (.CLK(clknet_leaf_130_clk),
    .D(_00579_),
    .Q(\regs[14][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14390_ (.CLK(clknet_leaf_2_clk),
    .D(_00580_),
    .Q(\regs[14][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14391_ (.CLK(clknet_leaf_105_clk),
    .D(_00581_),
    .Q(\regs[14][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14392_ (.CLK(clknet_leaf_127_clk),
    .D(_00582_),
    .Q(\regs[14][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14393_ (.CLK(clknet_leaf_2_clk),
    .D(_00583_),
    .Q(\regs[14][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14394_ (.CLK(clknet_leaf_106_clk),
    .D(_00584_),
    .Q(\regs[14][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14395_ (.CLK(clknet_leaf_104_clk),
    .D(_00585_),
    .Q(\regs[14][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14396_ (.CLK(clknet_leaf_98_clk),
    .D(_00586_),
    .Q(\regs[14][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14397_ (.CLK(clknet_leaf_104_clk),
    .D(_00587_),
    .Q(\regs[14][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14398_ (.CLK(clknet_leaf_90_clk),
    .D(_00588_),
    .Q(\regs[14][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14399_ (.CLK(clknet_leaf_99_clk),
    .D(_00589_),
    .Q(\regs[14][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14400_ (.CLK(clknet_leaf_107_clk),
    .D(_00590_),
    .Q(\regs[14][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14401_ (.CLK(clknet_leaf_99_clk),
    .D(_00591_),
    .Q(\regs[14][16] ));
 sky130_fd_sc_hd__dfxtp_1 _14402_ (.CLK(clknet_leaf_100_clk),
    .D(_00592_),
    .Q(\regs[14][17] ));
 sky130_fd_sc_hd__dfxtp_1 _14403_ (.CLK(clknet_leaf_100_clk),
    .D(_00593_),
    .Q(\regs[14][18] ));
 sky130_fd_sc_hd__dfxtp_1 _14404_ (.CLK(clknet_leaf_99_clk),
    .D(_00594_),
    .Q(\regs[14][19] ));
 sky130_fd_sc_hd__dfxtp_1 _14405_ (.CLK(clknet_leaf_9_clk),
    .D(_00595_),
    .Q(\regs[14][20] ));
 sky130_fd_sc_hd__dfxtp_1 _14406_ (.CLK(clknet_leaf_81_clk),
    .D(_00596_),
    .Q(\regs[14][21] ));
 sky130_fd_sc_hd__dfxtp_1 _14407_ (.CLK(clknet_leaf_65_clk),
    .D(_00597_),
    .Q(\regs[14][22] ));
 sky130_fd_sc_hd__dfxtp_1 _14408_ (.CLK(clknet_leaf_27_clk),
    .D(_00598_),
    .Q(\regs[14][23] ));
 sky130_fd_sc_hd__dfxtp_1 _14409_ (.CLK(clknet_leaf_20_clk),
    .D(_00599_),
    .Q(\regs[14][24] ));
 sky130_fd_sc_hd__dfxtp_1 _14410_ (.CLK(clknet_leaf_10_clk),
    .D(_00600_),
    .Q(\regs[14][25] ));
 sky130_fd_sc_hd__dfxtp_1 _14411_ (.CLK(clknet_leaf_70_clk),
    .D(_00601_),
    .Q(\regs[14][26] ));
 sky130_fd_sc_hd__dfxtp_1 _14412_ (.CLK(clknet_leaf_65_clk),
    .D(_00602_),
    .Q(\regs[14][27] ));
 sky130_fd_sc_hd__dfxtp_1 _14413_ (.CLK(clknet_leaf_10_clk),
    .D(_00603_),
    .Q(\regs[14][28] ));
 sky130_fd_sc_hd__dfxtp_1 _14414_ (.CLK(clknet_leaf_71_clk),
    .D(_00604_),
    .Q(\regs[14][29] ));
 sky130_fd_sc_hd__dfxtp_1 _14415_ (.CLK(clknet_leaf_115_clk),
    .D(_00605_),
    .Q(\regs[14][30] ));
 sky130_fd_sc_hd__dfxtp_1 _14416_ (.CLK(clknet_leaf_74_clk),
    .D(_00606_),
    .Q(\regs[14][31] ));
 sky130_fd_sc_hd__dfxtp_1 _14417_ (.CLK(clknet_leaf_118_clk),
    .D(_00607_),
    .Q(\regs[16][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14418_ (.CLK(clknet_leaf_132_clk),
    .D(_00608_),
    .Q(\regs[16][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14419_ (.CLK(clknet_leaf_132_clk),
    .D(_00609_),
    .Q(\regs[16][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14420_ (.CLK(clknet_leaf_2_clk),
    .D(_00610_),
    .Q(\regs[16][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14421_ (.CLK(clknet_leaf_122_clk),
    .D(_00611_),
    .Q(\regs[16][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14422_ (.CLK(clknet_leaf_4_clk),
    .D(_00612_),
    .Q(\regs[16][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14423_ (.CLK(clknet_leaf_107_clk),
    .D(_00613_),
    .Q(\regs[16][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14424_ (.CLK(clknet_leaf_124_clk),
    .D(_00614_),
    .Q(\regs[16][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14425_ (.CLK(clknet_leaf_4_clk),
    .D(_00615_),
    .Q(\regs[16][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14426_ (.CLK(clknet_leaf_124_clk),
    .D(_00616_),
    .Q(\regs[16][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14427_ (.CLK(clknet_leaf_75_clk),
    .D(_00617_),
    .Q(\regs[16][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14428_ (.CLK(clknet_leaf_87_clk),
    .D(_00618_),
    .Q(\regs[16][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14429_ (.CLK(clknet_leaf_88_clk),
    .D(_00619_),
    .Q(\regs[16][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14430_ (.CLK(clknet_leaf_86_clk),
    .D(_00620_),
    .Q(\regs[16][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14431_ (.CLK(clknet_leaf_85_clk),
    .D(_00621_),
    .Q(\regs[16][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14432_ (.CLK(clknet_leaf_112_clk),
    .D(_00622_),
    .Q(\regs[16][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14433_ (.CLK(clknet_leaf_82_clk),
    .D(_00623_),
    .Q(\regs[16][16] ));
 sky130_fd_sc_hd__dfxtp_1 _14434_ (.CLK(clknet_leaf_81_clk),
    .D(_00624_),
    .Q(\regs[16][17] ));
 sky130_fd_sc_hd__dfxtp_1 _14435_ (.CLK(clknet_leaf_76_clk),
    .D(_00625_),
    .Q(\regs[16][18] ));
 sky130_fd_sc_hd__dfxtp_1 _14436_ (.CLK(clknet_leaf_84_clk),
    .D(_00626_),
    .Q(\regs[16][19] ));
 sky130_fd_sc_hd__dfxtp_1 _14437_ (.CLK(clknet_leaf_26_clk),
    .D(_00627_),
    .Q(\regs[16][20] ));
 sky130_fd_sc_hd__dfxtp_1 _14438_ (.CLK(clknet_leaf_20_clk),
    .D(_00628_),
    .Q(\regs[16][21] ));
 sky130_fd_sc_hd__dfxtp_1 _14439_ (.CLK(clknet_leaf_55_clk),
    .D(_00629_),
    .Q(\regs[16][22] ));
 sky130_fd_sc_hd__dfxtp_1 _14440_ (.CLK(clknet_leaf_25_clk),
    .D(_00630_),
    .Q(\regs[16][23] ));
 sky130_fd_sc_hd__dfxtp_1 _14441_ (.CLK(clknet_leaf_23_clk),
    .D(_00631_),
    .Q(\regs[16][24] ));
 sky130_fd_sc_hd__dfxtp_1 _14442_ (.CLK(clknet_leaf_21_clk),
    .D(_00632_),
    .Q(\regs[16][25] ));
 sky130_fd_sc_hd__dfxtp_1 _14443_ (.CLK(clknet_leaf_53_clk),
    .D(_00633_),
    .Q(\regs[16][26] ));
 sky130_fd_sc_hd__dfxtp_1 _14444_ (.CLK(clknet_leaf_56_clk),
    .D(_00634_),
    .Q(\regs[16][27] ));
 sky130_fd_sc_hd__dfxtp_1 _14445_ (.CLK(clknet_leaf_26_clk),
    .D(_00635_),
    .Q(\regs[16][28] ));
 sky130_fd_sc_hd__dfxtp_1 _14446_ (.CLK(clknet_leaf_23_clk),
    .D(_00636_),
    .Q(\regs[16][29] ));
 sky130_fd_sc_hd__dfxtp_1 _14447_ (.CLK(clknet_leaf_55_clk),
    .D(_00637_),
    .Q(\regs[16][30] ));
 sky130_fd_sc_hd__dfxtp_1 _14448_ (.CLK(clknet_leaf_71_clk),
    .D(_00638_),
    .Q(\regs[16][31] ));
 sky130_fd_sc_hd__dfxtp_1 _14449_ (.CLK(clknet_leaf_125_clk),
    .D(_00639_),
    .Q(\regs[11][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14450_ (.CLK(clknet_leaf_133_clk),
    .D(_00640_),
    .Q(\regs[11][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14451_ (.CLK(clknet_leaf_128_clk),
    .D(_00641_),
    .Q(\regs[11][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14452_ (.CLK(clknet_leaf_135_clk),
    .D(_00642_),
    .Q(\regs[11][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14453_ (.CLK(clknet_leaf_128_clk),
    .D(_00643_),
    .Q(\regs[11][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14454_ (.CLK(clknet_leaf_2_clk),
    .D(_00644_),
    .Q(\regs[11][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14455_ (.CLK(clknet_leaf_105_clk),
    .D(_00645_),
    .Q(\regs[11][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14456_ (.CLK(clknet_leaf_126_clk),
    .D(_00646_),
    .Q(\regs[11][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14457_ (.CLK(clknet_leaf_135_clk),
    .D(_00647_),
    .Q(\regs[11][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14458_ (.CLK(clknet_leaf_105_clk),
    .D(_00648_),
    .Q(\regs[11][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14459_ (.CLK(clknet_leaf_103_clk),
    .D(_00649_),
    .Q(\regs[11][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14460_ (.CLK(clknet_leaf_98_clk),
    .D(_00650_),
    .Q(\regs[11][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14461_ (.CLK(clknet_leaf_102_clk),
    .D(_00651_),
    .Q(\regs[11][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14462_ (.CLK(clknet_leaf_101_clk),
    .D(_00652_),
    .Q(\regs[11][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14463_ (.CLK(clknet_leaf_97_clk),
    .D(_00653_),
    .Q(\regs[11][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14464_ (.CLK(clknet_leaf_104_clk),
    .D(_00654_),
    .Q(\regs[11][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14465_ (.CLK(clknet_leaf_97_clk),
    .D(_00655_),
    .Q(\regs[11][16] ));
 sky130_fd_sc_hd__dfxtp_1 _14466_ (.CLK(clknet_leaf_103_clk),
    .D(_00656_),
    .Q(\regs[11][17] ));
 sky130_fd_sc_hd__dfxtp_1 _14467_ (.CLK(clknet_leaf_101_clk),
    .D(_00657_),
    .Q(\regs[11][18] ));
 sky130_fd_sc_hd__dfxtp_1 _14468_ (.CLK(clknet_leaf_103_clk),
    .D(_00658_),
    .Q(\regs[11][19] ));
 sky130_fd_sc_hd__dfxtp_1 _14469_ (.CLK(clknet_leaf_6_clk),
    .D(_00659_),
    .Q(\regs[11][20] ));
 sky130_fd_sc_hd__dfxtp_1 _14470_ (.CLK(clknet_leaf_65_clk),
    .D(_00660_),
    .Q(\regs[11][21] ));
 sky130_fd_sc_hd__dfxtp_1 _14471_ (.CLK(clknet_leaf_66_clk),
    .D(_00661_),
    .Q(\regs[11][22] ));
 sky130_fd_sc_hd__dfxtp_1 _14472_ (.CLK(clknet_leaf_28_clk),
    .D(_00662_),
    .Q(\regs[11][23] ));
 sky130_fd_sc_hd__dfxtp_1 _14473_ (.CLK(clknet_leaf_20_clk),
    .D(_00663_),
    .Q(\regs[11][24] ));
 sky130_fd_sc_hd__dfxtp_1 _14474_ (.CLK(clknet_leaf_7_clk),
    .D(_00664_),
    .Q(\regs[11][25] ));
 sky130_fd_sc_hd__dfxtp_1 _14475_ (.CLK(clknet_leaf_66_clk),
    .D(_00665_),
    .Q(\regs[11][26] ));
 sky130_fd_sc_hd__dfxtp_1 _14476_ (.CLK(clknet_leaf_70_clk),
    .D(_00666_),
    .Q(\regs[11][27] ));
 sky130_fd_sc_hd__dfxtp_1 _14477_ (.CLK(clknet_leaf_7_clk),
    .D(_00667_),
    .Q(\regs[11][28] ));
 sky130_fd_sc_hd__dfxtp_1 _14478_ (.CLK(clknet_leaf_21_clk),
    .D(_00668_),
    .Q(\regs[11][29] ));
 sky130_fd_sc_hd__dfxtp_1 _14479_ (.CLK(clknet_leaf_114_clk),
    .D(_00669_),
    .Q(\regs[11][30] ));
 sky130_fd_sc_hd__dfxtp_1 _14480_ (.CLK(clknet_leaf_115_clk),
    .D(_00670_),
    .Q(\regs[11][31] ));
 sky130_fd_sc_hd__dfxtp_1 _14481_ (.CLK(clknet_leaf_120_clk),
    .D(_00671_),
    .Q(\regs[31][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14482_ (.CLK(clknet_leaf_14_clk),
    .D(_00672_),
    .Q(\regs[31][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14483_ (.CLK(clknet_leaf_121_clk),
    .D(_00673_),
    .Q(\regs[31][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14484_ (.CLK(clknet_leaf_3_clk),
    .D(_00674_),
    .Q(\regs[31][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14485_ (.CLK(clknet_leaf_122_clk),
    .D(_00675_),
    .Q(\regs[31][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14486_ (.CLK(clknet_leaf_13_clk),
    .D(_00676_),
    .Q(\regs[31][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14487_ (.CLK(clknet_leaf_108_clk),
    .D(_00677_),
    .Q(\regs[31][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14488_ (.CLK(clknet_leaf_123_clk),
    .D(_00678_),
    .Q(\regs[31][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14489_ (.CLK(clknet_leaf_3_clk),
    .D(_00679_),
    .Q(\regs[31][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14490_ (.CLK(clknet_leaf_118_clk),
    .D(_00680_),
    .Q(\regs[31][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14491_ (.CLK(clknet_leaf_111_clk),
    .D(_00681_),
    .Q(\regs[31][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14492_ (.CLK(clknet_leaf_89_clk),
    .D(_00682_),
    .Q(\regs[31][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14493_ (.CLK(clknet_leaf_89_clk),
    .D(_00683_),
    .Q(\regs[31][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14494_ (.CLK(clknet_leaf_89_clk),
    .D(_00684_),
    .Q(\regs[31][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14495_ (.CLK(clknet_leaf_79_clk),
    .D(_00685_),
    .Q(\regs[31][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14496_ (.CLK(clknet_leaf_113_clk),
    .D(_00686_),
    .Q(\regs[31][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14497_ (.CLK(clknet_leaf_89_clk),
    .D(_00687_),
    .Q(\regs[31][16] ));
 sky130_fd_sc_hd__dfxtp_1 _14498_ (.CLK(clknet_leaf_77_clk),
    .D(_00688_),
    .Q(\regs[31][17] ));
 sky130_fd_sc_hd__dfxtp_1 _14499_ (.CLK(clknet_leaf_78_clk),
    .D(_00689_),
    .Q(\regs[31][18] ));
 sky130_fd_sc_hd__dfxtp_1 _14500_ (.CLK(clknet_leaf_83_clk),
    .D(_00690_),
    .Q(\regs[31][19] ));
 sky130_fd_sc_hd__dfxtp_1 _14501_ (.CLK(clknet_leaf_12_clk),
    .D(_00691_),
    .Q(\regs[31][20] ));
 sky130_fd_sc_hd__dfxtp_1 _14502_ (.CLK(clknet_leaf_17_clk),
    .D(_00692_),
    .Q(\regs[31][21] ));
 sky130_fd_sc_hd__dfxtp_1 _14503_ (.CLK(clknet_leaf_73_clk),
    .D(_00693_),
    .Q(\regs[31][22] ));
 sky130_fd_sc_hd__dfxtp_1 _14504_ (.CLK(clknet_leaf_11_clk),
    .D(_00694_),
    .Q(\regs[31][23] ));
 sky130_fd_sc_hd__dfxtp_1 _14505_ (.CLK(clknet_leaf_17_clk),
    .D(_00695_),
    .Q(\regs[31][24] ));
 sky130_fd_sc_hd__dfxtp_1 _14506_ (.CLK(clknet_leaf_16_clk),
    .D(_00696_),
    .Q(\regs[31][25] ));
 sky130_fd_sc_hd__dfxtp_1 _14507_ (.CLK(clknet_leaf_19_clk),
    .D(_00697_),
    .Q(\regs[31][26] ));
 sky130_fd_sc_hd__dfxtp_1 _14508_ (.CLK(clknet_leaf_116_clk),
    .D(_00698_),
    .Q(\regs[31][27] ));
 sky130_fd_sc_hd__dfxtp_1 _14509_ (.CLK(clknet_leaf_10_clk),
    .D(_00699_),
    .Q(\regs[31][28] ));
 sky130_fd_sc_hd__dfxtp_1 _14510_ (.CLK(clknet_leaf_20_clk),
    .D(_00700_),
    .Q(\regs[31][29] ));
 sky130_fd_sc_hd__dfxtp_1 _14511_ (.CLK(clknet_leaf_115_clk),
    .D(_00701_),
    .Q(\regs[31][30] ));
 sky130_fd_sc_hd__dfxtp_1 _14512_ (.CLK(clknet_leaf_115_clk),
    .D(_00702_),
    .Q(\regs[31][31] ));
 sky130_fd_sc_hd__dfxtp_1 _14513_ (.CLK(clknet_leaf_15_clk),
    .D(_00703_),
    .Q(\regs[29][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14514_ (.CLK(clknet_leaf_15_clk),
    .D(_00704_),
    .Q(\regs[29][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14515_ (.CLK(clknet_leaf_121_clk),
    .D(_00705_),
    .Q(\regs[29][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14516_ (.CLK(clknet_leaf_3_clk),
    .D(_00706_),
    .Q(\regs[29][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14517_ (.CLK(clknet_leaf_122_clk),
    .D(_00707_),
    .Q(\regs[29][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14518_ (.CLK(clknet_leaf_13_clk),
    .D(_00708_),
    .Q(\regs[29][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14519_ (.CLK(clknet_leaf_108_clk),
    .D(_00709_),
    .Q(\regs[29][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14520_ (.CLK(clknet_leaf_123_clk),
    .D(_00710_),
    .Q(\regs[29][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14521_ (.CLK(clknet_leaf_3_clk),
    .D(_00711_),
    .Q(\regs[29][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14522_ (.CLK(clknet_leaf_114_clk),
    .D(_00712_),
    .Q(\regs[29][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14523_ (.CLK(clknet_leaf_111_clk),
    .D(_00713_),
    .Q(\regs[29][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14524_ (.CLK(clknet_leaf_89_clk),
    .D(_00714_),
    .Q(\regs[29][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14525_ (.CLK(clknet_leaf_90_clk),
    .D(_00715_),
    .Q(\regs[29][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14526_ (.CLK(clknet_leaf_89_clk),
    .D(_00716_),
    .Q(\regs[29][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14527_ (.CLK(clknet_leaf_82_clk),
    .D(_00717_),
    .Q(\regs[29][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14528_ (.CLK(clknet_leaf_113_clk),
    .D(_00718_),
    .Q(\regs[29][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14529_ (.CLK(clknet_leaf_90_clk),
    .D(_00719_),
    .Q(\regs[29][16] ));
 sky130_fd_sc_hd__dfxtp_1 _14530_ (.CLK(clknet_leaf_76_clk),
    .D(_00720_),
    .Q(\regs[29][17] ));
 sky130_fd_sc_hd__dfxtp_1 _14531_ (.CLK(clknet_leaf_112_clk),
    .D(_00721_),
    .Q(\regs[29][18] ));
 sky130_fd_sc_hd__dfxtp_1 _14532_ (.CLK(clknet_leaf_79_clk),
    .D(_00722_),
    .Q(\regs[29][19] ));
 sky130_fd_sc_hd__dfxtp_1 _14533_ (.CLK(clknet_leaf_11_clk),
    .D(_00723_),
    .Q(\regs[29][20] ));
 sky130_fd_sc_hd__dfxtp_1 _14534_ (.CLK(clknet_leaf_19_clk),
    .D(_00724_),
    .Q(\regs[29][21] ));
 sky130_fd_sc_hd__dfxtp_1 _14535_ (.CLK(clknet_leaf_116_clk),
    .D(_00725_),
    .Q(\regs[29][22] ));
 sky130_fd_sc_hd__dfxtp_1 _14536_ (.CLK(clknet_leaf_16_clk),
    .D(_00726_),
    .Q(\regs[29][23] ));
 sky130_fd_sc_hd__dfxtp_1 _14537_ (.CLK(clknet_leaf_21_clk),
    .D(_00727_),
    .Q(\regs[29][24] ));
 sky130_fd_sc_hd__dfxtp_1 _14538_ (.CLK(clknet_leaf_16_clk),
    .D(_00728_),
    .Q(\regs[29][25] ));
 sky130_fd_sc_hd__dfxtp_1 _14539_ (.CLK(clknet_leaf_19_clk),
    .D(_00729_),
    .Q(\regs[29][26] ));
 sky130_fd_sc_hd__dfxtp_1 _14540_ (.CLK(clknet_leaf_116_clk),
    .D(_00730_),
    .Q(\regs[29][27] ));
 sky130_fd_sc_hd__dfxtp_1 _14541_ (.CLK(clknet_leaf_11_clk),
    .D(_00731_),
    .Q(\regs[29][28] ));
 sky130_fd_sc_hd__dfxtp_1 _14542_ (.CLK(clknet_leaf_19_clk),
    .D(_00732_),
    .Q(\regs[29][29] ));
 sky130_fd_sc_hd__dfxtp_1 _14543_ (.CLK(clknet_leaf_116_clk),
    .D(_00733_),
    .Q(\regs[29][30] ));
 sky130_fd_sc_hd__dfxtp_1 _14544_ (.CLK(clknet_leaf_115_clk),
    .D(_00734_),
    .Q(\regs[29][31] ));
 sky130_fd_sc_hd__dfxtp_1 _14545_ (.CLK(clknet_leaf_122_clk),
    .D(_00735_),
    .Q(\regs[3][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14546_ (.CLK(clknet_leaf_134_clk),
    .D(_00736_),
    .Q(\regs[3][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14547_ (.CLK(clknet_leaf_129_clk),
    .D(_00737_),
    .Q(\regs[3][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14548_ (.CLK(clknet_leaf_0_clk),
    .D(_00738_),
    .Q(\regs[3][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14549_ (.CLK(clknet_leaf_131_clk),
    .D(_00739_),
    .Q(\regs[3][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14550_ (.CLK(clknet_leaf_5_clk),
    .D(_00740_),
    .Q(\regs[3][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14551_ (.CLK(clknet_leaf_126_clk),
    .D(_00741_),
    .Q(\regs[3][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14552_ (.CLK(clknet_leaf_127_clk),
    .D(_00742_),
    .Q(\regs[3][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14553_ (.CLK(clknet_leaf_0_clk),
    .D(_00743_),
    .Q(\regs[3][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14554_ (.CLK(clknet_leaf_106_clk),
    .D(_00744_),
    .Q(\regs[3][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14555_ (.CLK(clknet_leaf_101_clk),
    .D(_00745_),
    .Q(\regs[3][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14556_ (.CLK(clknet_leaf_95_clk),
    .D(_00746_),
    .Q(\regs[3][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14557_ (.CLK(clknet_leaf_102_clk),
    .D(_00747_),
    .Q(\regs[3][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14558_ (.CLK(clknet_leaf_92_clk),
    .D(_00748_),
    .Q(\regs[3][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14559_ (.CLK(clknet_leaf_93_clk),
    .D(_00749_),
    .Q(\regs[3][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14560_ (.CLK(clknet_leaf_109_clk),
    .D(_00750_),
    .Q(\regs[3][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14561_ (.CLK(clknet_leaf_94_clk),
    .D(_00751_),
    .Q(\regs[3][16] ));
 sky130_fd_sc_hd__dfxtp_1 _14562_ (.CLK(clknet_leaf_100_clk),
    .D(_00752_),
    .Q(\regs[3][17] ));
 sky130_fd_sc_hd__dfxtp_1 _14563_ (.CLK(clknet_leaf_110_clk),
    .D(_00753_),
    .Q(\regs[3][18] ));
 sky130_fd_sc_hd__dfxtp_1 _14564_ (.CLK(clknet_leaf_92_clk),
    .D(_00754_),
    .Q(\regs[3][19] ));
 sky130_fd_sc_hd__dfxtp_1 _14565_ (.CLK(clknet_leaf_8_clk),
    .D(_00755_),
    .Q(\regs[3][20] ));
 sky130_fd_sc_hd__dfxtp_1 _14566_ (.CLK(clknet_leaf_63_clk),
    .D(_00756_),
    .Q(\regs[3][21] ));
 sky130_fd_sc_hd__dfxtp_1 _14567_ (.CLK(clknet_leaf_64_clk),
    .D(_00757_),
    .Q(\regs[3][22] ));
 sky130_fd_sc_hd__dfxtp_1 _14568_ (.CLK(clknet_leaf_30_clk),
    .D(_00758_),
    .Q(\regs[3][23] ));
 sky130_fd_sc_hd__dfxtp_1 _14569_ (.CLK(clknet_leaf_26_clk),
    .D(_00759_),
    .Q(\regs[3][24] ));
 sky130_fd_sc_hd__dfxtp_1 _14570_ (.CLK(clknet_leaf_9_clk),
    .D(_00760_),
    .Q(\regs[3][25] ));
 sky130_fd_sc_hd__dfxtp_1 _14571_ (.CLK(clknet_leaf_71_clk),
    .D(_00761_),
    .Q(\regs[3][26] ));
 sky130_fd_sc_hd__dfxtp_1 _14572_ (.CLK(clknet_leaf_64_clk),
    .D(_00762_),
    .Q(\regs[3][27] ));
 sky130_fd_sc_hd__dfxtp_1 _14573_ (.CLK(clknet_leaf_29_clk),
    .D(_00763_),
    .Q(\regs[3][28] ));
 sky130_fd_sc_hd__dfxtp_1 _14574_ (.CLK(clknet_leaf_71_clk),
    .D(_00764_),
    .Q(\regs[3][29] ));
 sky130_fd_sc_hd__dfxtp_1 _14575_ (.CLK(clknet_leaf_73_clk),
    .D(_00765_),
    .Q(\regs[3][30] ));
 sky130_fd_sc_hd__dfxtp_1 _14576_ (.CLK(clknet_leaf_74_clk),
    .D(_00766_),
    .Q(\regs[3][31] ));
 sky130_fd_sc_hd__dfxtp_1 _14577_ (.CLK(clknet_leaf_119_clk),
    .D(_00767_),
    .Q(\regs[19][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14578_ (.CLK(clknet_leaf_132_clk),
    .D(_00768_),
    .Q(\regs[19][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14579_ (.CLK(clknet_leaf_132_clk),
    .D(_00769_),
    .Q(\regs[19][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14580_ (.CLK(clknet_leaf_4_clk),
    .D(_00770_),
    .Q(\regs[19][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14581_ (.CLK(clknet_leaf_121_clk),
    .D(_00771_),
    .Q(\regs[19][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14582_ (.CLK(clknet_leaf_4_clk),
    .D(_00772_),
    .Q(\regs[19][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14583_ (.CLK(clknet_leaf_108_clk),
    .D(_00773_),
    .Q(\regs[19][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14584_ (.CLK(clknet_leaf_122_clk),
    .D(_00774_),
    .Q(\regs[19][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14585_ (.CLK(clknet_leaf_4_clk),
    .D(_00775_),
    .Q(\regs[19][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14586_ (.CLK(clknet_leaf_124_clk),
    .D(_00776_),
    .Q(\regs[19][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14587_ (.CLK(clknet_leaf_70_clk),
    .D(_00777_),
    .Q(\regs[19][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14588_ (.CLK(clknet_leaf_86_clk),
    .D(_00778_),
    .Q(\regs[19][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14589_ (.CLK(clknet_leaf_87_clk),
    .D(_00779_),
    .Q(\regs[19][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14590_ (.CLK(clknet_leaf_85_clk),
    .D(_00780_),
    .Q(\regs[19][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14591_ (.CLK(clknet_leaf_85_clk),
    .D(_00781_),
    .Q(\regs[19][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14592_ (.CLK(clknet_leaf_112_clk),
    .D(_00782_),
    .Q(\regs[19][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14593_ (.CLK(clknet_leaf_83_clk),
    .D(_00783_),
    .Q(\regs[19][16] ));
 sky130_fd_sc_hd__dfxtp_1 _14594_ (.CLK(clknet_leaf_81_clk),
    .D(_00784_),
    .Q(\regs[19][17] ));
 sky130_fd_sc_hd__dfxtp_1 _14595_ (.CLK(clknet_leaf_76_clk),
    .D(_00785_),
    .Q(\regs[19][18] ));
 sky130_fd_sc_hd__dfxtp_1 _14596_ (.CLK(clknet_leaf_84_clk),
    .D(_00786_),
    .Q(\regs[19][19] ));
 sky130_fd_sc_hd__dfxtp_1 _14597_ (.CLK(clknet_leaf_27_clk),
    .D(_00787_),
    .Q(\regs[19][20] ));
 sky130_fd_sc_hd__dfxtp_1 _14598_ (.CLK(clknet_leaf_20_clk),
    .D(_00788_),
    .Q(\regs[19][21] ));
 sky130_fd_sc_hd__dfxtp_1 _14599_ (.CLK(clknet_leaf_53_clk),
    .D(_00789_),
    .Q(\regs[19][22] ));
 sky130_fd_sc_hd__dfxtp_1 _14600_ (.CLK(clknet_leaf_25_clk),
    .D(_00790_),
    .Q(\regs[19][23] ));
 sky130_fd_sc_hd__dfxtp_1 _14601_ (.CLK(clknet_leaf_24_clk),
    .D(_00791_),
    .Q(\regs[19][24] ));
 sky130_fd_sc_hd__dfxtp_1 _14602_ (.CLK(clknet_leaf_16_clk),
    .D(_00792_),
    .Q(\regs[19][25] ));
 sky130_fd_sc_hd__dfxtp_1 _14603_ (.CLK(clknet_leaf_53_clk),
    .D(_00793_),
    .Q(\regs[19][26] ));
 sky130_fd_sc_hd__dfxtp_1 _14604_ (.CLK(clknet_leaf_56_clk),
    .D(_00794_),
    .Q(\regs[19][27] ));
 sky130_fd_sc_hd__dfxtp_1 _14605_ (.CLK(clknet_leaf_26_clk),
    .D(_00795_),
    .Q(\regs[19][28] ));
 sky130_fd_sc_hd__dfxtp_1 _14606_ (.CLK(clknet_leaf_23_clk),
    .D(_00796_),
    .Q(\regs[19][29] ));
 sky130_fd_sc_hd__dfxtp_1 _14607_ (.CLK(clknet_leaf_55_clk),
    .D(_00797_),
    .Q(\regs[19][30] ));
 sky130_fd_sc_hd__dfxtp_1 _14608_ (.CLK(clknet_leaf_71_clk),
    .D(_00798_),
    .Q(\regs[19][31] ));
 sky130_fd_sc_hd__dfxtp_1 _14609_ (.CLK(clknet_leaf_125_clk),
    .D(_00799_),
    .Q(\regs[4][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14610_ (.CLK(clknet_leaf_130_clk),
    .D(_00800_),
    .Q(\regs[4][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14611_ (.CLK(clknet_leaf_129_clk),
    .D(_00801_),
    .Q(\regs[4][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14612_ (.CLK(clknet_leaf_2_clk),
    .D(_00802_),
    .Q(\regs[4][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14613_ (.CLK(clknet_leaf_130_clk),
    .D(_00803_),
    .Q(\regs[4][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14614_ (.CLK(clknet_leaf_2_clk),
    .D(_00804_),
    .Q(\regs[4][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14615_ (.CLK(clknet_leaf_105_clk),
    .D(_00805_),
    .Q(\regs[4][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14616_ (.CLK(clknet_leaf_126_clk),
    .D(_00806_),
    .Q(\regs[4][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14617_ (.CLK(clknet_leaf_1_clk),
    .D(_00807_),
    .Q(\regs[4][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14618_ (.CLK(clknet_leaf_106_clk),
    .D(_00808_),
    .Q(\regs[4][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14619_ (.CLK(clknet_leaf_100_clk),
    .D(_00809_),
    .Q(\regs[4][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14620_ (.CLK(clknet_leaf_96_clk),
    .D(_00810_),
    .Q(\regs[4][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14621_ (.CLK(clknet_leaf_98_clk),
    .D(_00811_),
    .Q(\regs[4][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14622_ (.CLK(clknet_leaf_92_clk),
    .D(_00812_),
    .Q(\regs[4][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14623_ (.CLK(clknet_leaf_95_clk),
    .D(_00813_),
    .Q(\regs[4][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14624_ (.CLK(clknet_leaf_109_clk),
    .D(_00814_),
    .Q(\regs[4][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14625_ (.CLK(clknet_leaf_91_clk),
    .D(_00815_),
    .Q(\regs[4][16] ));
 sky130_fd_sc_hd__dfxtp_1 _14626_ (.CLK(clknet_leaf_100_clk),
    .D(_00816_),
    .Q(\regs[4][17] ));
 sky130_fd_sc_hd__dfxtp_1 _14627_ (.CLK(clknet_leaf_100_clk),
    .D(_00817_),
    .Q(\regs[4][18] ));
 sky130_fd_sc_hd__dfxtp_1 _14628_ (.CLK(clknet_leaf_92_clk),
    .D(_00818_),
    .Q(\regs[4][19] ));
 sky130_fd_sc_hd__dfxtp_1 _14629_ (.CLK(clknet_leaf_7_clk),
    .D(_00819_),
    .Q(\regs[4][20] ));
 sky130_fd_sc_hd__dfxtp_1 _14630_ (.CLK(clknet_leaf_64_clk),
    .D(_00820_),
    .Q(\regs[4][21] ));
 sky130_fd_sc_hd__dfxtp_1 _14631_ (.CLK(clknet_leaf_64_clk),
    .D(_00821_),
    .Q(\regs[4][22] ));
 sky130_fd_sc_hd__dfxtp_1 _14632_ (.CLK(clknet_leaf_28_clk),
    .D(_00822_),
    .Q(\regs[4][23] ));
 sky130_fd_sc_hd__dfxtp_1 _14633_ (.CLK(clknet_leaf_22_clk),
    .D(_00823_),
    .Q(\regs[4][24] ));
 sky130_fd_sc_hd__dfxtp_1 _14634_ (.CLK(clknet_leaf_9_clk),
    .D(_00824_),
    .Q(\regs[4][25] ));
 sky130_fd_sc_hd__dfxtp_1 _14635_ (.CLK(clknet_leaf_69_clk),
    .D(_00825_),
    .Q(\regs[4][26] ));
 sky130_fd_sc_hd__dfxtp_1 _14636_ (.CLK(clknet_leaf_66_clk),
    .D(_00826_),
    .Q(\regs[4][27] ));
 sky130_fd_sc_hd__dfxtp_1 _14637_ (.CLK(clknet_leaf_29_clk),
    .D(_00827_),
    .Q(\regs[4][28] ));
 sky130_fd_sc_hd__dfxtp_1 _14638_ (.CLK(clknet_leaf_20_clk),
    .D(_00828_),
    .Q(\regs[4][29] ));
 sky130_fd_sc_hd__dfxtp_1 _14639_ (.CLK(clknet_leaf_73_clk),
    .D(_00829_),
    .Q(\regs[4][30] ));
 sky130_fd_sc_hd__dfxtp_1 _14640_ (.CLK(clknet_leaf_74_clk),
    .D(_00830_),
    .Q(\regs[4][31] ));
 sky130_fd_sc_hd__dfrtp_2 _14641_ (.CLK(clknet_leaf_51_clk),
    .D(_00831_),
    .RESET_B(_00072_),
    .Q(\PC[1] ));
 sky130_fd_sc_hd__dfxtp_1 _14642_ (.CLK(clknet_leaf_125_clk),
    .D(_00832_),
    .Q(\regs[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14643_ (.CLK(clknet_leaf_129_clk),
    .D(_00833_),
    .Q(\regs[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14644_ (.CLK(clknet_leaf_129_clk),
    .D(_00834_),
    .Q(\regs[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14645_ (.CLK(clknet_leaf_135_clk),
    .D(_00835_),
    .Q(\regs[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14646_ (.CLK(clknet_leaf_130_clk),
    .D(_00836_),
    .Q(\regs[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14647_ (.CLK(clknet_leaf_0_clk),
    .D(_00837_),
    .Q(\regs[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14648_ (.CLK(clknet_leaf_105_clk),
    .D(_00838_),
    .Q(\regs[0][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14649_ (.CLK(clknet_leaf_127_clk),
    .D(_00839_),
    .Q(\regs[0][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14650_ (.CLK(clknet_leaf_1_clk),
    .D(_00840_),
    .Q(\regs[0][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14651_ (.CLK(clknet_leaf_107_clk),
    .D(_00841_),
    .Q(\regs[0][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14652_ (.CLK(clknet_leaf_101_clk),
    .D(_00842_),
    .Q(\regs[0][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14653_ (.CLK(clknet_leaf_95_clk),
    .D(_00843_),
    .Q(\regs[0][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14654_ (.CLK(clknet_leaf_102_clk),
    .D(_00844_),
    .Q(\regs[0][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14655_ (.CLK(clknet_leaf_92_clk),
    .D(_00845_),
    .Q(\regs[0][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14656_ (.CLK(clknet_leaf_95_clk),
    .D(_00846_),
    .Q(\regs[0][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14657_ (.CLK(clknet_leaf_110_clk),
    .D(_00847_),
    .Q(\regs[0][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14658_ (.CLK(clknet_leaf_93_clk),
    .D(_00848_),
    .Q(\regs[0][16] ));
 sky130_fd_sc_hd__dfxtp_1 _14659_ (.CLK(clknet_leaf_90_clk),
    .D(_00849_),
    .Q(\regs[0][17] ));
 sky130_fd_sc_hd__dfxtp_1 _14660_ (.CLK(clknet_leaf_111_clk),
    .D(_00850_),
    .Q(\regs[0][18] ));
 sky130_fd_sc_hd__dfxtp_1 _14661_ (.CLK(clknet_leaf_85_clk),
    .D(_00851_),
    .Q(\regs[0][19] ));
 sky130_fd_sc_hd__dfxtp_1 _14662_ (.CLK(clknet_leaf_8_clk),
    .D(_00852_),
    .Q(\regs[0][20] ));
 sky130_fd_sc_hd__dfxtp_1 _14663_ (.CLK(clknet_leaf_63_clk),
    .D(_00853_),
    .Q(\regs[0][21] ));
 sky130_fd_sc_hd__dfxtp_1 _14664_ (.CLK(clknet_leaf_63_clk),
    .D(_00854_),
    .Q(\regs[0][22] ));
 sky130_fd_sc_hd__dfxtp_1 _14665_ (.CLK(clknet_leaf_28_clk),
    .D(_00855_),
    .Q(\regs[0][23] ));
 sky130_fd_sc_hd__dfxtp_1 _14666_ (.CLK(clknet_leaf_26_clk),
    .D(_00856_),
    .Q(\regs[0][24] ));
 sky130_fd_sc_hd__dfxtp_1 _14667_ (.CLK(clknet_leaf_8_clk),
    .D(_00857_),
    .Q(\regs[0][25] ));
 sky130_fd_sc_hd__dfxtp_1 _14668_ (.CLK(clknet_leaf_69_clk),
    .D(_00858_),
    .Q(\regs[0][26] ));
 sky130_fd_sc_hd__dfxtp_1 _14669_ (.CLK(clknet_leaf_64_clk),
    .D(_00859_),
    .Q(\regs[0][27] ));
 sky130_fd_sc_hd__dfxtp_1 _14670_ (.CLK(clknet_leaf_29_clk),
    .D(_00860_),
    .Q(\regs[0][28] ));
 sky130_fd_sc_hd__dfxtp_1 _14671_ (.CLK(clknet_leaf_71_clk),
    .D(_00861_),
    .Q(\regs[0][29] ));
 sky130_fd_sc_hd__dfxtp_1 _14672_ (.CLK(clknet_leaf_74_clk),
    .D(_00862_),
    .Q(\regs[0][30] ));
 sky130_fd_sc_hd__dfxtp_1 _14673_ (.CLK(clknet_leaf_75_clk),
    .D(_00863_),
    .Q(\regs[0][31] ));
 sky130_fd_sc_hd__dfxtp_1 _14674_ (.CLK(clknet_leaf_119_clk),
    .D(_00864_),
    .Q(\regs[18][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14675_ (.CLK(clknet_leaf_132_clk),
    .D(_00865_),
    .Q(\regs[18][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14676_ (.CLK(clknet_leaf_132_clk),
    .D(_00866_),
    .Q(\regs[18][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14677_ (.CLK(clknet_leaf_4_clk),
    .D(_00867_),
    .Q(\regs[18][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14678_ (.CLK(clknet_leaf_122_clk),
    .D(_00868_),
    .Q(\regs[18][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14679_ (.CLK(clknet_leaf_4_clk),
    .D(_00869_),
    .Q(\regs[18][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14680_ (.CLK(clknet_leaf_108_clk),
    .D(_00870_),
    .Q(\regs[18][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14681_ (.CLK(clknet_leaf_122_clk),
    .D(_00871_),
    .Q(\regs[18][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14682_ (.CLK(clknet_leaf_4_clk),
    .D(_00872_),
    .Q(\regs[18][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14683_ (.CLK(clknet_leaf_124_clk),
    .D(_00873_),
    .Q(\regs[18][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14684_ (.CLK(clknet_leaf_70_clk),
    .D(_00874_),
    .Q(\regs[18][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14685_ (.CLK(clknet_leaf_88_clk),
    .D(_00875_),
    .Q(\regs[18][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14686_ (.CLK(clknet_leaf_88_clk),
    .D(_00876_),
    .Q(\regs[18][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14687_ (.CLK(clknet_leaf_86_clk),
    .D(_00877_),
    .Q(\regs[18][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14688_ (.CLK(clknet_leaf_83_clk),
    .D(_00878_),
    .Q(\regs[18][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14689_ (.CLK(clknet_leaf_112_clk),
    .D(_00879_),
    .Q(\regs[18][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14690_ (.CLK(clknet_leaf_82_clk),
    .D(_00880_),
    .Q(\regs[18][16] ));
 sky130_fd_sc_hd__dfxtp_1 _14691_ (.CLK(clknet_leaf_75_clk),
    .D(_00881_),
    .Q(\regs[18][17] ));
 sky130_fd_sc_hd__dfxtp_1 _14692_ (.CLK(clknet_leaf_74_clk),
    .D(_00882_),
    .Q(\regs[18][18] ));
 sky130_fd_sc_hd__dfxtp_1 _14693_ (.CLK(clknet_leaf_83_clk),
    .D(_00883_),
    .Q(\regs[18][19] ));
 sky130_fd_sc_hd__dfxtp_1 _14694_ (.CLK(clknet_leaf_27_clk),
    .D(_00884_),
    .Q(\regs[18][20] ));
 sky130_fd_sc_hd__dfxtp_1 _14695_ (.CLK(clknet_leaf_20_clk),
    .D(_00885_),
    .Q(\regs[18][21] ));
 sky130_fd_sc_hd__dfxtp_1 _14696_ (.CLK(clknet_leaf_53_clk),
    .D(_00886_),
    .Q(\regs[18][22] ));
 sky130_fd_sc_hd__dfxtp_1 _14697_ (.CLK(clknet_leaf_25_clk),
    .D(_00887_),
    .Q(\regs[18][23] ));
 sky130_fd_sc_hd__dfxtp_1 _14698_ (.CLK(clknet_leaf_24_clk),
    .D(_00888_),
    .Q(\regs[18][24] ));
 sky130_fd_sc_hd__dfxtp_1 _14699_ (.CLK(clknet_leaf_21_clk),
    .D(_00889_),
    .Q(\regs[18][25] ));
 sky130_fd_sc_hd__dfxtp_1 _14700_ (.CLK(clknet_leaf_54_clk),
    .D(_00890_),
    .Q(\regs[18][26] ));
 sky130_fd_sc_hd__dfxtp_1 _14701_ (.CLK(clknet_leaf_56_clk),
    .D(_00891_),
    .Q(\regs[18][27] ));
 sky130_fd_sc_hd__dfxtp_1 _14702_ (.CLK(clknet_leaf_27_clk),
    .D(_00892_),
    .Q(\regs[18][28] ));
 sky130_fd_sc_hd__dfxtp_1 _14703_ (.CLK(clknet_leaf_23_clk),
    .D(_00893_),
    .Q(\regs[18][29] ));
 sky130_fd_sc_hd__dfxtp_1 _14704_ (.CLK(clknet_leaf_55_clk),
    .D(_00894_),
    .Q(\regs[18][30] ));
 sky130_fd_sc_hd__dfxtp_1 _14705_ (.CLK(clknet_leaf_71_clk),
    .D(_00895_),
    .Q(\regs[18][31] ));
 sky130_fd_sc_hd__dfxtp_1 _14706_ (.CLK(clknet_leaf_125_clk),
    .D(_00896_),
    .Q(\regs[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14707_ (.CLK(clknet_leaf_134_clk),
    .D(_00897_),
    .Q(\regs[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14708_ (.CLK(clknet_leaf_129_clk),
    .D(_00898_),
    .Q(\regs[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14709_ (.CLK(clknet_leaf_0_clk),
    .D(_00899_),
    .Q(\regs[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14710_ (.CLK(clknet_leaf_130_clk),
    .D(_00900_),
    .Q(\regs[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14711_ (.CLK(clknet_leaf_5_clk),
    .D(_00901_),
    .Q(\regs[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14712_ (.CLK(clknet_leaf_105_clk),
    .D(_00902_),
    .Q(\regs[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14713_ (.CLK(clknet_leaf_127_clk),
    .D(_00903_),
    .Q(\regs[1][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14714_ (.CLK(clknet_leaf_0_clk),
    .D(_00904_),
    .Q(\regs[1][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14715_ (.CLK(clknet_leaf_106_clk),
    .D(_00905_),
    .Q(\regs[1][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14716_ (.CLK(clknet_leaf_101_clk),
    .D(_00906_),
    .Q(\regs[1][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14717_ (.CLK(clknet_leaf_95_clk),
    .D(_00907_),
    .Q(\regs[1][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14718_ (.CLK(clknet_leaf_102_clk),
    .D(_00908_),
    .Q(\regs[1][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14719_ (.CLK(clknet_leaf_92_clk),
    .D(_00909_),
    .Q(\regs[1][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14720_ (.CLK(clknet_leaf_93_clk),
    .D(_00910_),
    .Q(\regs[1][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14721_ (.CLK(clknet_leaf_110_clk),
    .D(_00911_),
    .Q(\regs[1][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14722_ (.CLK(clknet_leaf_93_clk),
    .D(_00912_),
    .Q(\regs[1][16] ));
 sky130_fd_sc_hd__dfxtp_1 _14723_ (.CLK(clknet_leaf_100_clk),
    .D(_00913_),
    .Q(\regs[1][17] ));
 sky130_fd_sc_hd__dfxtp_1 _14724_ (.CLK(clknet_leaf_111_clk),
    .D(_00914_),
    .Q(\regs[1][18] ));
 sky130_fd_sc_hd__dfxtp_1 _14725_ (.CLK(clknet_leaf_93_clk),
    .D(_00915_),
    .Q(\regs[1][19] ));
 sky130_fd_sc_hd__dfxtp_1 _14726_ (.CLK(clknet_leaf_8_clk),
    .D(_00916_),
    .Q(\regs[1][20] ));
 sky130_fd_sc_hd__dfxtp_1 _14727_ (.CLK(clknet_leaf_63_clk),
    .D(_00917_),
    .Q(\regs[1][21] ));
 sky130_fd_sc_hd__dfxtp_1 _14728_ (.CLK(clknet_leaf_63_clk),
    .D(_00918_),
    .Q(\regs[1][22] ));
 sky130_fd_sc_hd__dfxtp_1 _14729_ (.CLK(clknet_leaf_30_clk),
    .D(_00919_),
    .Q(\regs[1][23] ));
 sky130_fd_sc_hd__dfxtp_1 _14730_ (.CLK(clknet_leaf_26_clk),
    .D(_00920_),
    .Q(\regs[1][24] ));
 sky130_fd_sc_hd__dfxtp_1 _14731_ (.CLK(clknet_leaf_9_clk),
    .D(_00921_),
    .Q(\regs[1][25] ));
 sky130_fd_sc_hd__dfxtp_1 _14732_ (.CLK(clknet_leaf_68_clk),
    .D(_00922_),
    .Q(\regs[1][26] ));
 sky130_fd_sc_hd__dfxtp_1 _14733_ (.CLK(clknet_leaf_64_clk),
    .D(_00923_),
    .Q(\regs[1][27] ));
 sky130_fd_sc_hd__dfxtp_1 _14734_ (.CLK(clknet_leaf_29_clk),
    .D(_00924_),
    .Q(\regs[1][28] ));
 sky130_fd_sc_hd__dfxtp_1 _14735_ (.CLK(clknet_leaf_71_clk),
    .D(_00925_),
    .Q(\regs[1][29] ));
 sky130_fd_sc_hd__dfxtp_1 _14736_ (.CLK(clknet_leaf_72_clk),
    .D(_00926_),
    .Q(\regs[1][30] ));
 sky130_fd_sc_hd__dfxtp_1 _14737_ (.CLK(clknet_leaf_75_clk),
    .D(_00927_),
    .Q(\regs[1][31] ));
 sky130_fd_sc_hd__dfxtp_1 _14738_ (.CLK(clknet_leaf_118_clk),
    .D(_00928_),
    .Q(\regs[20][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14739_ (.CLK(clknet_leaf_132_clk),
    .D(_00929_),
    .Q(\regs[20][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14740_ (.CLK(clknet_leaf_131_clk),
    .D(_00930_),
    .Q(\regs[20][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14741_ (.CLK(clknet_leaf_4_clk),
    .D(_00931_),
    .Q(\regs[20][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14742_ (.CLK(clknet_leaf_122_clk),
    .D(_00932_),
    .Q(\regs[20][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14743_ (.CLK(clknet_leaf_4_clk),
    .D(_00933_),
    .Q(\regs[20][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14744_ (.CLK(clknet_leaf_107_clk),
    .D(_00934_),
    .Q(\regs[20][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14745_ (.CLK(clknet_leaf_125_clk),
    .D(_00935_),
    .Q(\regs[20][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14746_ (.CLK(clknet_leaf_4_clk),
    .D(_00936_),
    .Q(\regs[20][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14747_ (.CLK(clknet_leaf_108_clk),
    .D(_00937_),
    .Q(\regs[20][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14748_ (.CLK(clknet_leaf_75_clk),
    .D(_00938_),
    .Q(\regs[20][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14749_ (.CLK(clknet_leaf_87_clk),
    .D(_00939_),
    .Q(\regs[20][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14750_ (.CLK(clknet_leaf_87_clk),
    .D(_00940_),
    .Q(\regs[20][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14751_ (.CLK(clknet_leaf_86_clk),
    .D(_00941_),
    .Q(\regs[20][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14752_ (.CLK(clknet_leaf_85_clk),
    .D(_00942_),
    .Q(\regs[20][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14753_ (.CLK(clknet_leaf_112_clk),
    .D(_00943_),
    .Q(\regs[20][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14754_ (.CLK(clknet_leaf_84_clk),
    .D(_00944_),
    .Q(\regs[20][16] ));
 sky130_fd_sc_hd__dfxtp_1 _14755_ (.CLK(clknet_leaf_80_clk),
    .D(_00945_),
    .Q(\regs[20][17] ));
 sky130_fd_sc_hd__dfxtp_1 _14756_ (.CLK(clknet_leaf_80_clk),
    .D(_00946_),
    .Q(\regs[20][18] ));
 sky130_fd_sc_hd__dfxtp_1 _14757_ (.CLK(clknet_leaf_84_clk),
    .D(_00947_),
    .Q(\regs[20][19] ));
 sky130_fd_sc_hd__dfxtp_1 _14758_ (.CLK(clknet_leaf_27_clk),
    .D(_00948_),
    .Q(\regs[20][20] ));
 sky130_fd_sc_hd__dfxtp_1 _14759_ (.CLK(clknet_leaf_20_clk),
    .D(_00949_),
    .Q(\regs[20][21] ));
 sky130_fd_sc_hd__dfxtp_1 _14760_ (.CLK(clknet_leaf_55_clk),
    .D(_00950_),
    .Q(\regs[20][22] ));
 sky130_fd_sc_hd__dfxtp_1 _14761_ (.CLK(clknet_leaf_25_clk),
    .D(_00951_),
    .Q(\regs[20][23] ));
 sky130_fd_sc_hd__dfxtp_1 _14762_ (.CLK(clknet_leaf_20_clk),
    .D(_00952_),
    .Q(\regs[20][24] ));
 sky130_fd_sc_hd__dfxtp_1 _14763_ (.CLK(clknet_leaf_21_clk),
    .D(_00953_),
    .Q(\regs[20][25] ));
 sky130_fd_sc_hd__dfxtp_1 _14764_ (.CLK(clknet_leaf_54_clk),
    .D(_00954_),
    .Q(\regs[20][26] ));
 sky130_fd_sc_hd__dfxtp_1 _14765_ (.CLK(clknet_leaf_56_clk),
    .D(_00955_),
    .Q(\regs[20][27] ));
 sky130_fd_sc_hd__dfxtp_1 _14766_ (.CLK(clknet_leaf_27_clk),
    .D(_00956_),
    .Q(\regs[20][28] ));
 sky130_fd_sc_hd__dfxtp_1 _14767_ (.CLK(clknet_leaf_22_clk),
    .D(_00957_),
    .Q(\regs[20][29] ));
 sky130_fd_sc_hd__dfxtp_1 _14768_ (.CLK(clknet_leaf_72_clk),
    .D(_00958_),
    .Q(\regs[20][30] ));
 sky130_fd_sc_hd__dfxtp_1 _14769_ (.CLK(clknet_leaf_70_clk),
    .D(_00959_),
    .Q(\regs[20][31] ));
 sky130_fd_sc_hd__dfxtp_1 _14770_ (.CLK(clknet_leaf_119_clk),
    .D(_00960_),
    .Q(\regs[21][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14771_ (.CLK(clknet_leaf_132_clk),
    .D(_00961_),
    .Q(\regs[21][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14772_ (.CLK(clknet_leaf_131_clk),
    .D(_00962_),
    .Q(\regs[21][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14773_ (.CLK(clknet_leaf_5_clk),
    .D(_00963_),
    .Q(\regs[21][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14774_ (.CLK(clknet_leaf_122_clk),
    .D(_00964_),
    .Q(\regs[21][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14775_ (.CLK(clknet_leaf_6_clk),
    .D(_00965_),
    .Q(\regs[21][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14776_ (.CLK(clknet_leaf_107_clk),
    .D(_00966_),
    .Q(\regs[21][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14777_ (.CLK(clknet_leaf_125_clk),
    .D(_00967_),
    .Q(\regs[21][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14778_ (.CLK(clknet_leaf_6_clk),
    .D(_00968_),
    .Q(\regs[21][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14779_ (.CLK(clknet_leaf_124_clk),
    .D(_00969_),
    .Q(\regs[21][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14780_ (.CLK(clknet_leaf_75_clk),
    .D(_00970_),
    .Q(\regs[21][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14781_ (.CLK(clknet_leaf_87_clk),
    .D(_00971_),
    .Q(\regs[21][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14782_ (.CLK(clknet_leaf_87_clk),
    .D(_00972_),
    .Q(\regs[21][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14783_ (.CLK(clknet_leaf_85_clk),
    .D(_00973_),
    .Q(\regs[21][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14784_ (.CLK(clknet_leaf_85_clk),
    .D(_00974_),
    .Q(\regs[21][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14785_ (.CLK(clknet_leaf_110_clk),
    .D(_00975_),
    .Q(\regs[21][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14786_ (.CLK(clknet_leaf_85_clk),
    .D(_00976_),
    .Q(\regs[21][16] ));
 sky130_fd_sc_hd__dfxtp_1 _14787_ (.CLK(clknet_leaf_80_clk),
    .D(_00977_),
    .Q(\regs[21][17] ));
 sky130_fd_sc_hd__dfxtp_1 _14788_ (.CLK(clknet_leaf_80_clk),
    .D(_00978_),
    .Q(\regs[21][18] ));
 sky130_fd_sc_hd__dfxtp_1 _14789_ (.CLK(clknet_leaf_84_clk),
    .D(_00979_),
    .Q(\regs[21][19] ));
 sky130_fd_sc_hd__dfxtp_1 _14790_ (.CLK(clknet_leaf_28_clk),
    .D(_00980_),
    .Q(\regs[21][20] ));
 sky130_fd_sc_hd__dfxtp_1 _14791_ (.CLK(clknet_leaf_20_clk),
    .D(_00981_),
    .Q(\regs[21][21] ));
 sky130_fd_sc_hd__dfxtp_1 _14792_ (.CLK(clknet_leaf_55_clk),
    .D(_00982_),
    .Q(\regs[21][22] ));
 sky130_fd_sc_hd__dfxtp_1 _14793_ (.CLK(clknet_leaf_25_clk),
    .D(_00983_),
    .Q(\regs[21][23] ));
 sky130_fd_sc_hd__dfxtp_1 _14794_ (.CLK(clknet_leaf_22_clk),
    .D(_00984_),
    .Q(\regs[21][24] ));
 sky130_fd_sc_hd__dfxtp_1 _14795_ (.CLK(clknet_leaf_21_clk),
    .D(_00985_),
    .Q(\regs[21][25] ));
 sky130_fd_sc_hd__dfxtp_1 _14796_ (.CLK(clknet_leaf_54_clk),
    .D(_00986_),
    .Q(\regs[21][26] ));
 sky130_fd_sc_hd__dfxtp_1 _14797_ (.CLK(clknet_leaf_55_clk),
    .D(_00987_),
    .Q(\regs[21][27] ));
 sky130_fd_sc_hd__dfxtp_1 _14798_ (.CLK(clknet_leaf_28_clk),
    .D(_00988_),
    .Q(\regs[21][28] ));
 sky130_fd_sc_hd__dfxtp_1 _14799_ (.CLK(clknet_leaf_23_clk),
    .D(_00989_),
    .Q(\regs[21][29] ));
 sky130_fd_sc_hd__dfxtp_1 _14800_ (.CLK(clknet_leaf_72_clk),
    .D(_00990_),
    .Q(\regs[21][30] ));
 sky130_fd_sc_hd__dfxtp_1 _14801_ (.CLK(clknet_leaf_70_clk),
    .D(_00991_),
    .Q(\regs[21][31] ));
 sky130_fd_sc_hd__dfxtp_1 _14802_ (.CLK(clknet_leaf_119_clk),
    .D(_00992_),
    .Q(\regs[22][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14803_ (.CLK(clknet_leaf_133_clk),
    .D(_00993_),
    .Q(\regs[22][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14804_ (.CLK(clknet_leaf_132_clk),
    .D(_00994_),
    .Q(\regs[22][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14805_ (.CLK(clknet_leaf_5_clk),
    .D(_00995_),
    .Q(\regs[22][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14806_ (.CLK(clknet_leaf_131_clk),
    .D(_00996_),
    .Q(\regs[22][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14807_ (.CLK(clknet_leaf_6_clk),
    .D(_00997_),
    .Q(\regs[22][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14808_ (.CLK(clknet_leaf_108_clk),
    .D(_00998_),
    .Q(\regs[22][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14809_ (.CLK(clknet_leaf_122_clk),
    .D(_00999_),
    .Q(\regs[22][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14810_ (.CLK(clknet_leaf_6_clk),
    .D(_01000_),
    .Q(\regs[22][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14811_ (.CLK(clknet_leaf_124_clk),
    .D(_01001_),
    .Q(\regs[22][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14812_ (.CLK(clknet_leaf_75_clk),
    .D(_01002_),
    .Q(\regs[22][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14813_ (.CLK(clknet_leaf_87_clk),
    .D(_01003_),
    .Q(\regs[22][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14814_ (.CLK(clknet_leaf_87_clk),
    .D(_01004_),
    .Q(\regs[22][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14815_ (.CLK(clknet_leaf_86_clk),
    .D(_01005_),
    .Q(\regs[22][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14816_ (.CLK(clknet_leaf_85_clk),
    .D(_01006_),
    .Q(\regs[22][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14817_ (.CLK(clknet_leaf_113_clk),
    .D(_01007_),
    .Q(\regs[22][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14818_ (.CLK(clknet_leaf_83_clk),
    .D(_01008_),
    .Q(\regs[22][16] ));
 sky130_fd_sc_hd__dfxtp_1 _14819_ (.CLK(clknet_leaf_76_clk),
    .D(_01009_),
    .Q(\regs[22][17] ));
 sky130_fd_sc_hd__dfxtp_1 _14820_ (.CLK(clknet_leaf_76_clk),
    .D(_01010_),
    .Q(\regs[22][18] ));
 sky130_fd_sc_hd__dfxtp_1 _14821_ (.CLK(clknet_leaf_84_clk),
    .D(_01011_),
    .Q(\regs[22][19] ));
 sky130_fd_sc_hd__dfxtp_1 _14822_ (.CLK(clknet_leaf_29_clk),
    .D(_01012_),
    .Q(\regs[22][20] ));
 sky130_fd_sc_hd__dfxtp_1 _14823_ (.CLK(clknet_leaf_22_clk),
    .D(_01013_),
    .Q(\regs[22][21] ));
 sky130_fd_sc_hd__dfxtp_1 _14824_ (.CLK(clknet_leaf_55_clk),
    .D(_01014_),
    .Q(\regs[22][22] ));
 sky130_fd_sc_hd__dfxtp_1 _14825_ (.CLK(clknet_leaf_28_clk),
    .D(_01015_),
    .Q(\regs[22][23] ));
 sky130_fd_sc_hd__dfxtp_1 _14826_ (.CLK(clknet_leaf_22_clk),
    .D(_01016_),
    .Q(\regs[22][24] ));
 sky130_fd_sc_hd__dfxtp_1 _14827_ (.CLK(clknet_leaf_26_clk),
    .D(_01017_),
    .Q(\regs[22][25] ));
 sky130_fd_sc_hd__dfxtp_1 _14828_ (.CLK(clknet_leaf_54_clk),
    .D(_01018_),
    .Q(\regs[22][26] ));
 sky130_fd_sc_hd__dfxtp_1 _14829_ (.CLK(clknet_leaf_55_clk),
    .D(_01019_),
    .Q(\regs[22][27] ));
 sky130_fd_sc_hd__dfxtp_1 _14830_ (.CLK(clknet_leaf_28_clk),
    .D(_01020_),
    .Q(\regs[22][28] ));
 sky130_fd_sc_hd__dfxtp_1 _14831_ (.CLK(clknet_leaf_22_clk),
    .D(_01021_),
    .Q(\regs[22][29] ));
 sky130_fd_sc_hd__dfxtp_1 _14832_ (.CLK(clknet_leaf_72_clk),
    .D(_01022_),
    .Q(\regs[22][30] ));
 sky130_fd_sc_hd__dfxtp_1 _14833_ (.CLK(clknet_leaf_70_clk),
    .D(_01023_),
    .Q(\regs[22][31] ));
 sky130_fd_sc_hd__dfxtp_1 _14834_ (.CLK(clknet_leaf_119_clk),
    .D(_01024_),
    .Q(\regs[23][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14835_ (.CLK(clknet_leaf_132_clk),
    .D(_01025_),
    .Q(\regs[23][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14836_ (.CLK(clknet_leaf_132_clk),
    .D(_01026_),
    .Q(\regs[23][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14837_ (.CLK(clknet_leaf_5_clk),
    .D(_01027_),
    .Q(\regs[23][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14838_ (.CLK(clknet_leaf_122_clk),
    .D(_01028_),
    .Q(\regs[23][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14839_ (.CLK(clknet_leaf_6_clk),
    .D(_01029_),
    .Q(\regs[23][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14840_ (.CLK(clknet_leaf_107_clk),
    .D(_01030_),
    .Q(\regs[23][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14841_ (.CLK(clknet_leaf_122_clk),
    .D(_01031_),
    .Q(\regs[23][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14842_ (.CLK(clknet_leaf_5_clk),
    .D(_01032_),
    .Q(\regs[23][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14843_ (.CLK(clknet_leaf_124_clk),
    .D(_01033_),
    .Q(\regs[23][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14844_ (.CLK(clknet_leaf_80_clk),
    .D(_01034_),
    .Q(\regs[23][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14845_ (.CLK(clknet_leaf_87_clk),
    .D(_01035_),
    .Q(\regs[23][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14846_ (.CLK(clknet_leaf_87_clk),
    .D(_01036_),
    .Q(\regs[23][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14847_ (.CLK(clknet_leaf_86_clk),
    .D(_01037_),
    .Q(\regs[23][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14848_ (.CLK(clknet_leaf_85_clk),
    .D(_01038_),
    .Q(\regs[23][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14849_ (.CLK(clknet_leaf_113_clk),
    .D(_01039_),
    .Q(\regs[23][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14850_ (.CLK(clknet_leaf_85_clk),
    .D(_01040_),
    .Q(\regs[23][16] ));
 sky130_fd_sc_hd__dfxtp_1 _14851_ (.CLK(clknet_leaf_80_clk),
    .D(_01041_),
    .Q(\regs[23][17] ));
 sky130_fd_sc_hd__dfxtp_1 _14852_ (.CLK(clknet_leaf_76_clk),
    .D(_01042_),
    .Q(\regs[23][18] ));
 sky130_fd_sc_hd__dfxtp_1 _14853_ (.CLK(clknet_leaf_84_clk),
    .D(_01043_),
    .Q(\regs[23][19] ));
 sky130_fd_sc_hd__dfxtp_1 _14854_ (.CLK(clknet_leaf_29_clk),
    .D(_01044_),
    .Q(\regs[23][20] ));
 sky130_fd_sc_hd__dfxtp_1 _14855_ (.CLK(clknet_leaf_20_clk),
    .D(_01045_),
    .Q(\regs[23][21] ));
 sky130_fd_sc_hd__dfxtp_1 _14856_ (.CLK(clknet_leaf_55_clk),
    .D(_01046_),
    .Q(\regs[23][22] ));
 sky130_fd_sc_hd__dfxtp_1 _14857_ (.CLK(clknet_leaf_28_clk),
    .D(_01047_),
    .Q(\regs[23][23] ));
 sky130_fd_sc_hd__dfxtp_1 _14858_ (.CLK(clknet_leaf_22_clk),
    .D(_01048_),
    .Q(\regs[23][24] ));
 sky130_fd_sc_hd__dfxtp_1 _14859_ (.CLK(clknet_leaf_26_clk),
    .D(_01049_),
    .Q(\regs[23][25] ));
 sky130_fd_sc_hd__dfxtp_1 _14860_ (.CLK(clknet_leaf_54_clk),
    .D(_01050_),
    .Q(\regs[23][26] ));
 sky130_fd_sc_hd__dfxtp_1 _14861_ (.CLK(clknet_leaf_55_clk),
    .D(_01051_),
    .Q(\regs[23][27] ));
 sky130_fd_sc_hd__dfxtp_1 _14862_ (.CLK(clknet_leaf_28_clk),
    .D(_01052_),
    .Q(\regs[23][28] ));
 sky130_fd_sc_hd__dfxtp_1 _14863_ (.CLK(clknet_leaf_23_clk),
    .D(_01053_),
    .Q(\regs[23][29] ));
 sky130_fd_sc_hd__dfxtp_1 _14864_ (.CLK(clknet_leaf_72_clk),
    .D(_01054_),
    .Q(\regs[23][30] ));
 sky130_fd_sc_hd__dfxtp_1 _14865_ (.CLK(clknet_leaf_71_clk),
    .D(_01055_),
    .Q(\regs[23][31] ));
 sky130_fd_sc_hd__dfxtp_1 _14866_ (.CLK(clknet_leaf_117_clk),
    .D(_01056_),
    .Q(\regs[24][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14867_ (.CLK(clknet_leaf_14_clk),
    .D(_01057_),
    .Q(\regs[24][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14868_ (.CLK(clknet_leaf_121_clk),
    .D(_01058_),
    .Q(\regs[24][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14869_ (.CLK(clknet_leaf_132_clk),
    .D(_01059_),
    .Q(\regs[24][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14870_ (.CLK(clknet_leaf_121_clk),
    .D(_01060_),
    .Q(\regs[24][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14871_ (.CLK(clknet_leaf_14_clk),
    .D(_01061_),
    .Q(\regs[24][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14872_ (.CLK(clknet_leaf_123_clk),
    .D(_01062_),
    .Q(\regs[24][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14873_ (.CLK(clknet_leaf_123_clk),
    .D(_01063_),
    .Q(\regs[24][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14874_ (.CLK(clknet_leaf_14_clk),
    .D(_01064_),
    .Q(\regs[24][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14875_ (.CLK(clknet_leaf_118_clk),
    .D(_01065_),
    .Q(\regs[24][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14876_ (.CLK(clknet_leaf_111_clk),
    .D(_01066_),
    .Q(\regs[24][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14877_ (.CLK(clknet_leaf_78_clk),
    .D(_01067_),
    .Q(\regs[24][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14878_ (.CLK(clknet_leaf_90_clk),
    .D(_01068_),
    .Q(\regs[24][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14879_ (.CLK(clknet_leaf_77_clk),
    .D(_01069_),
    .Q(\regs[24][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14880_ (.CLK(clknet_leaf_79_clk),
    .D(_01070_),
    .Q(\regs[24][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14881_ (.CLK(clknet_leaf_114_clk),
    .D(_01071_),
    .Q(\regs[24][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14882_ (.CLK(clknet_leaf_90_clk),
    .D(_01072_),
    .Q(\regs[24][16] ));
 sky130_fd_sc_hd__dfxtp_1 _14883_ (.CLK(clknet_leaf_77_clk),
    .D(_01073_),
    .Q(\regs[24][17] ));
 sky130_fd_sc_hd__dfxtp_1 _14884_ (.CLK(clknet_leaf_78_clk),
    .D(_01074_),
    .Q(\regs[24][18] ));
 sky130_fd_sc_hd__dfxtp_1 _14885_ (.CLK(clknet_leaf_80_clk),
    .D(_01075_),
    .Q(\regs[24][19] ));
 sky130_fd_sc_hd__dfxtp_1 _14886_ (.CLK(clknet_leaf_14_clk),
    .D(_01076_),
    .Q(\regs[24][20] ));
 sky130_fd_sc_hd__dfxtp_1 _14887_ (.CLK(clknet_leaf_17_clk),
    .D(_01077_),
    .Q(\regs[24][21] ));
 sky130_fd_sc_hd__dfxtp_1 _14888_ (.CLK(clknet_leaf_117_clk),
    .D(_01078_),
    .Q(\regs[24][22] ));
 sky130_fd_sc_hd__dfxtp_1 _14889_ (.CLK(clknet_leaf_11_clk),
    .D(_01079_),
    .Q(\regs[24][23] ));
 sky130_fd_sc_hd__dfxtp_1 _14890_ (.CLK(clknet_leaf_17_clk),
    .D(_01080_),
    .Q(\regs[24][24] ));
 sky130_fd_sc_hd__dfxtp_1 _14891_ (.CLK(clknet_leaf_15_clk),
    .D(_01081_),
    .Q(\regs[24][25] ));
 sky130_fd_sc_hd__dfxtp_1 _14892_ (.CLK(clknet_leaf_19_clk),
    .D(_01082_),
    .Q(\regs[24][26] ));
 sky130_fd_sc_hd__dfxtp_1 _14893_ (.CLK(clknet_leaf_117_clk),
    .D(_01083_),
    .Q(\regs[24][27] ));
 sky130_fd_sc_hd__dfxtp_1 _14894_ (.CLK(clknet_leaf_11_clk),
    .D(_01084_),
    .Q(\regs[24][28] ));
 sky130_fd_sc_hd__dfxtp_1 _14895_ (.CLK(clknet_leaf_15_clk),
    .D(_01085_),
    .Q(\regs[24][29] ));
 sky130_fd_sc_hd__dfxtp_1 _14896_ (.CLK(clknet_leaf_118_clk),
    .D(_01086_),
    .Q(\regs[24][30] ));
 sky130_fd_sc_hd__dfxtp_1 _14897_ (.CLK(clknet_leaf_117_clk),
    .D(_01087_),
    .Q(\regs[24][31] ));
 sky130_fd_sc_hd__dfxtp_1 _14898_ (.CLK(clknet_leaf_117_clk),
    .D(_01088_),
    .Q(\regs[25][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14899_ (.CLK(clknet_leaf_121_clk),
    .D(_01089_),
    .Q(\regs[25][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14900_ (.CLK(clknet_leaf_121_clk),
    .D(_01090_),
    .Q(\regs[25][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14901_ (.CLK(clknet_leaf_132_clk),
    .D(_01091_),
    .Q(\regs[25][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14902_ (.CLK(clknet_leaf_121_clk),
    .D(_01092_),
    .Q(\regs[25][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14903_ (.CLK(clknet_leaf_14_clk),
    .D(_01093_),
    .Q(\regs[25][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14904_ (.CLK(clknet_leaf_124_clk),
    .D(_01094_),
    .Q(\regs[25][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14905_ (.CLK(clknet_leaf_123_clk),
    .D(_01095_),
    .Q(\regs[25][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14906_ (.CLK(clknet_leaf_14_clk),
    .D(_01096_),
    .Q(\regs[25][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14907_ (.CLK(clknet_leaf_118_clk),
    .D(_01097_),
    .Q(\regs[25][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14908_ (.CLK(clknet_leaf_111_clk),
    .D(_01098_),
    .Q(\regs[25][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14909_ (.CLK(clknet_leaf_78_clk),
    .D(_01099_),
    .Q(\regs[25][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14910_ (.CLK(clknet_leaf_90_clk),
    .D(_01100_),
    .Q(\regs[25][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14911_ (.CLK(clknet_leaf_78_clk),
    .D(_01101_),
    .Q(\regs[25][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14912_ (.CLK(clknet_leaf_79_clk),
    .D(_01102_),
    .Q(\regs[25][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14913_ (.CLK(clknet_leaf_113_clk),
    .D(_01103_),
    .Q(\regs[25][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14914_ (.CLK(clknet_leaf_90_clk),
    .D(_01104_),
    .Q(\regs[25][16] ));
 sky130_fd_sc_hd__dfxtp_1 _14915_ (.CLK(clknet_leaf_77_clk),
    .D(_01105_),
    .Q(\regs[25][17] ));
 sky130_fd_sc_hd__dfxtp_1 _14916_ (.CLK(clknet_leaf_78_clk),
    .D(_01106_),
    .Q(\regs[25][18] ));
 sky130_fd_sc_hd__dfxtp_1 _14917_ (.CLK(clknet_leaf_79_clk),
    .D(_01107_),
    .Q(\regs[25][19] ));
 sky130_fd_sc_hd__dfxtp_1 _14918_ (.CLK(clknet_leaf_14_clk),
    .D(_01108_),
    .Q(\regs[25][20] ));
 sky130_fd_sc_hd__dfxtp_1 _14919_ (.CLK(clknet_leaf_17_clk),
    .D(_01109_),
    .Q(\regs[25][21] ));
 sky130_fd_sc_hd__dfxtp_1 _14920_ (.CLK(clknet_leaf_117_clk),
    .D(_01110_),
    .Q(\regs[25][22] ));
 sky130_fd_sc_hd__dfxtp_1 _14921_ (.CLK(clknet_leaf_16_clk),
    .D(_01111_),
    .Q(\regs[25][23] ));
 sky130_fd_sc_hd__dfxtp_1 _14922_ (.CLK(clknet_leaf_17_clk),
    .D(_01112_),
    .Q(\regs[25][24] ));
 sky130_fd_sc_hd__dfxtp_1 _14923_ (.CLK(clknet_leaf_15_clk),
    .D(_01113_),
    .Q(\regs[25][25] ));
 sky130_fd_sc_hd__dfxtp_1 _14924_ (.CLK(clknet_leaf_19_clk),
    .D(_01114_),
    .Q(\regs[25][26] ));
 sky130_fd_sc_hd__dfxtp_1 _14925_ (.CLK(clknet_leaf_117_clk),
    .D(_01115_),
    .Q(\regs[25][27] ));
 sky130_fd_sc_hd__dfxtp_1 _14926_ (.CLK(clknet_leaf_12_clk),
    .D(_01116_),
    .Q(\regs[25][28] ));
 sky130_fd_sc_hd__dfxtp_1 _14927_ (.CLK(clknet_leaf_18_clk),
    .D(_01117_),
    .Q(\regs[25][29] ));
 sky130_fd_sc_hd__dfxtp_1 _14928_ (.CLK(clknet_leaf_114_clk),
    .D(_01118_),
    .Q(\regs[25][30] ));
 sky130_fd_sc_hd__dfxtp_1 _14929_ (.CLK(clknet_leaf_117_clk),
    .D(_01119_),
    .Q(\regs[25][31] ));
 sky130_fd_sc_hd__dfxtp_1 _14930_ (.CLK(clknet_leaf_120_clk),
    .D(_01120_),
    .Q(\regs[26][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14931_ (.CLK(clknet_leaf_14_clk),
    .D(_01121_),
    .Q(\regs[26][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14932_ (.CLK(clknet_leaf_121_clk),
    .D(_01122_),
    .Q(\regs[26][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14933_ (.CLK(clknet_leaf_121_clk),
    .D(_01123_),
    .Q(\regs[26][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14934_ (.CLK(clknet_leaf_119_clk),
    .D(_01124_),
    .Q(\regs[26][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14935_ (.CLK(clknet_leaf_13_clk),
    .D(_01125_),
    .Q(\regs[26][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14936_ (.CLK(clknet_leaf_124_clk),
    .D(_01126_),
    .Q(\regs[26][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14937_ (.CLK(clknet_leaf_123_clk),
    .D(_01127_),
    .Q(\regs[26][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14938_ (.CLK(clknet_leaf_3_clk),
    .D(_01128_),
    .Q(\regs[26][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14939_ (.CLK(clknet_leaf_118_clk),
    .D(_01129_),
    .Q(\regs[26][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14940_ (.CLK(clknet_leaf_112_clk),
    .D(_01130_),
    .Q(\regs[26][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14941_ (.CLK(clknet_leaf_78_clk),
    .D(_01131_),
    .Q(\regs[26][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14942_ (.CLK(clknet_leaf_111_clk),
    .D(_01132_),
    .Q(\regs[26][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14943_ (.CLK(clknet_leaf_78_clk),
    .D(_01133_),
    .Q(\regs[26][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14944_ (.CLK(clknet_leaf_80_clk),
    .D(_01134_),
    .Q(\regs[26][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14945_ (.CLK(clknet_leaf_113_clk),
    .D(_01135_),
    .Q(\regs[26][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14946_ (.CLK(clknet_leaf_78_clk),
    .D(_01136_),
    .Q(\regs[26][16] ));
 sky130_fd_sc_hd__dfxtp_1 _14947_ (.CLK(clknet_leaf_74_clk),
    .D(_01137_),
    .Q(\regs[26][17] ));
 sky130_fd_sc_hd__dfxtp_1 _14948_ (.CLK(clknet_leaf_78_clk),
    .D(_01138_),
    .Q(\regs[26][18] ));
 sky130_fd_sc_hd__dfxtp_1 _14949_ (.CLK(clknet_leaf_79_clk),
    .D(_01139_),
    .Q(\regs[26][19] ));
 sky130_fd_sc_hd__dfxtp_1 _14950_ (.CLK(clknet_leaf_13_clk),
    .D(_01140_),
    .Q(\regs[26][20] ));
 sky130_fd_sc_hd__dfxtp_1 _14951_ (.CLK(clknet_leaf_18_clk),
    .D(_01141_),
    .Q(\regs[26][21] ));
 sky130_fd_sc_hd__dfxtp_1 _14952_ (.CLK(clknet_leaf_117_clk),
    .D(_01142_),
    .Q(\regs[26][22] ));
 sky130_fd_sc_hd__dfxtp_1 _14953_ (.CLK(clknet_leaf_15_clk),
    .D(_01143_),
    .Q(\regs[26][23] ));
 sky130_fd_sc_hd__dfxtp_1 _14954_ (.CLK(clknet_leaf_17_clk),
    .D(_01144_),
    .Q(\regs[26][24] ));
 sky130_fd_sc_hd__dfxtp_1 _14955_ (.CLK(clknet_leaf_15_clk),
    .D(_01145_),
    .Q(\regs[26][25] ));
 sky130_fd_sc_hd__dfxtp_1 _14956_ (.CLK(clknet_leaf_18_clk),
    .D(_01146_),
    .Q(\regs[26][26] ));
 sky130_fd_sc_hd__dfxtp_1 _14957_ (.CLK(clknet_leaf_117_clk),
    .D(_01147_),
    .Q(\regs[26][27] ));
 sky130_fd_sc_hd__dfxtp_1 _14958_ (.CLK(clknet_leaf_12_clk),
    .D(_01148_),
    .Q(\regs[26][28] ));
 sky130_fd_sc_hd__dfxtp_1 _14959_ (.CLK(clknet_leaf_18_clk),
    .D(_01149_),
    .Q(\regs[26][29] ));
 sky130_fd_sc_hd__dfxtp_1 _14960_ (.CLK(clknet_leaf_115_clk),
    .D(_01150_),
    .Q(\regs[26][30] ));
 sky130_fd_sc_hd__dfxtp_1 _14961_ (.CLK(clknet_leaf_117_clk),
    .D(_01151_),
    .Q(\regs[26][31] ));
 sky130_fd_sc_hd__dfxtp_1 _14962_ (.CLK(clknet_leaf_125_clk),
    .D(_01152_),
    .Q(\regs[6][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14963_ (.CLK(clknet_leaf_134_clk),
    .D(_01153_),
    .Q(\regs[6][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14964_ (.CLK(clknet_leaf_129_clk),
    .D(_01154_),
    .Q(\regs[6][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14965_ (.CLK(clknet_leaf_0_clk),
    .D(_01155_),
    .Q(\regs[6][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14966_ (.CLK(clknet_leaf_131_clk),
    .D(_01156_),
    .Q(\regs[6][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14967_ (.CLK(clknet_leaf_1_clk),
    .D(_01157_),
    .Q(\regs[6][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14968_ (.CLK(clknet_leaf_105_clk),
    .D(_01158_),
    .Q(\regs[6][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14969_ (.CLK(clknet_leaf_127_clk),
    .D(_01159_),
    .Q(\regs[6][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14970_ (.CLK(clknet_leaf_1_clk),
    .D(_01160_),
    .Q(\regs[6][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14971_ (.CLK(clknet_leaf_125_clk),
    .D(_01161_),
    .Q(\regs[6][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14972_ (.CLK(clknet_leaf_110_clk),
    .D(_01162_),
    .Q(\regs[6][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14973_ (.CLK(clknet_leaf_96_clk),
    .D(_01163_),
    .Q(\regs[6][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14974_ (.CLK(clknet_leaf_98_clk),
    .D(_01164_),
    .Q(\regs[6][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14975_ (.CLK(clknet_leaf_92_clk),
    .D(_01165_),
    .Q(\regs[6][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14976_ (.CLK(clknet_leaf_91_clk),
    .D(_01166_),
    .Q(\regs[6][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14977_ (.CLK(clknet_leaf_109_clk),
    .D(_01167_),
    .Q(\regs[6][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14978_ (.CLK(clknet_leaf_91_clk),
    .D(_01168_),
    .Q(\regs[6][16] ));
 sky130_fd_sc_hd__dfxtp_1 _14979_ (.CLK(clknet_leaf_100_clk),
    .D(_01169_),
    .Q(\regs[6][17] ));
 sky130_fd_sc_hd__dfxtp_1 _14980_ (.CLK(clknet_leaf_111_clk),
    .D(_01170_),
    .Q(\regs[6][18] ));
 sky130_fd_sc_hd__dfxtp_1 _14981_ (.CLK(clknet_leaf_91_clk),
    .D(_01171_),
    .Q(\regs[6][19] ));
 sky130_fd_sc_hd__dfxtp_1 _14982_ (.CLK(clknet_leaf_8_clk),
    .D(_01172_),
    .Q(\regs[6][20] ));
 sky130_fd_sc_hd__dfxtp_1 _14983_ (.CLK(clknet_leaf_64_clk),
    .D(_01173_),
    .Q(\regs[6][21] ));
 sky130_fd_sc_hd__dfxtp_1 _14984_ (.CLK(clknet_leaf_64_clk),
    .D(_01174_),
    .Q(\regs[6][22] ));
 sky130_fd_sc_hd__dfxtp_1 _14985_ (.CLK(clknet_leaf_28_clk),
    .D(_01175_),
    .Q(\regs[6][23] ));
 sky130_fd_sc_hd__dfxtp_1 _14986_ (.CLK(clknet_leaf_25_clk),
    .D(_01176_),
    .Q(\regs[6][24] ));
 sky130_fd_sc_hd__dfxtp_1 _14987_ (.CLK(clknet_leaf_9_clk),
    .D(_01177_),
    .Q(\regs[6][25] ));
 sky130_fd_sc_hd__dfxtp_1 _14988_ (.CLK(clknet_leaf_68_clk),
    .D(_01178_),
    .Q(\regs[6][26] ));
 sky130_fd_sc_hd__dfxtp_1 _14989_ (.CLK(clknet_leaf_66_clk),
    .D(_01179_),
    .Q(\regs[6][27] ));
 sky130_fd_sc_hd__dfxtp_1 _14990_ (.CLK(clknet_leaf_29_clk),
    .D(_01180_),
    .Q(\regs[6][28] ));
 sky130_fd_sc_hd__dfxtp_1 _14991_ (.CLK(clknet_leaf_71_clk),
    .D(_01181_),
    .Q(\regs[6][29] ));
 sky130_fd_sc_hd__dfxtp_1 _14992_ (.CLK(clknet_leaf_116_clk),
    .D(_01182_),
    .Q(\regs[6][30] ));
 sky130_fd_sc_hd__dfxtp_1 _14993_ (.CLK(clknet_leaf_74_clk),
    .D(_01183_),
    .Q(\regs[6][31] ));
 sky130_fd_sc_hd__dfxtp_1 _14994_ (.CLK(clknet_leaf_120_clk),
    .D(_01184_),
    .Q(\regs[27][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14995_ (.CLK(clknet_leaf_14_clk),
    .D(_01185_),
    .Q(\regs[27][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14996_ (.CLK(clknet_leaf_121_clk),
    .D(_01186_),
    .Q(\regs[27][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14997_ (.CLK(clknet_leaf_3_clk),
    .D(_01187_),
    .Q(\regs[27][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14998_ (.CLK(clknet_leaf_120_clk),
    .D(_01188_),
    .Q(\regs[27][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14999_ (.CLK(clknet_leaf_13_clk),
    .D(_01189_),
    .Q(\regs[27][5] ));
 sky130_fd_sc_hd__dfxtp_1 _15000_ (.CLK(clknet_leaf_123_clk),
    .D(_01190_),
    .Q(\regs[27][6] ));
 sky130_fd_sc_hd__dfxtp_1 _15001_ (.CLK(clknet_leaf_123_clk),
    .D(_01191_),
    .Q(\regs[27][7] ));
 sky130_fd_sc_hd__dfxtp_1 _15002_ (.CLK(clknet_leaf_13_clk),
    .D(_01192_),
    .Q(\regs[27][8] ));
 sky130_fd_sc_hd__dfxtp_1 _15003_ (.CLK(clknet_leaf_118_clk),
    .D(_01193_),
    .Q(\regs[27][9] ));
 sky130_fd_sc_hd__dfxtp_1 _15004_ (.CLK(clknet_leaf_111_clk),
    .D(_01194_),
    .Q(\regs[27][10] ));
 sky130_fd_sc_hd__dfxtp_1 _15005_ (.CLK(clknet_leaf_78_clk),
    .D(_01195_),
    .Q(\regs[27][11] ));
 sky130_fd_sc_hd__dfxtp_1 _15006_ (.CLK(clknet_leaf_111_clk),
    .D(_01196_),
    .Q(\regs[27][12] ));
 sky130_fd_sc_hd__dfxtp_1 _15007_ (.CLK(clknet_leaf_78_clk),
    .D(_01197_),
    .Q(\regs[27][13] ));
 sky130_fd_sc_hd__dfxtp_1 _15008_ (.CLK(clknet_leaf_80_clk),
    .D(_01198_),
    .Q(\regs[27][14] ));
 sky130_fd_sc_hd__dfxtp_1 _15009_ (.CLK(clknet_leaf_114_clk),
    .D(_01199_),
    .Q(\regs[27][15] ));
 sky130_fd_sc_hd__dfxtp_1 _15010_ (.CLK(clknet_leaf_78_clk),
    .D(_01200_),
    .Q(\regs[27][16] ));
 sky130_fd_sc_hd__dfxtp_1 _15011_ (.CLK(clknet_leaf_77_clk),
    .D(_01201_),
    .Q(\regs[27][17] ));
 sky130_fd_sc_hd__dfxtp_1 _15012_ (.CLK(clknet_leaf_111_clk),
    .D(_01202_),
    .Q(\regs[27][18] ));
 sky130_fd_sc_hd__dfxtp_1 _15013_ (.CLK(clknet_leaf_79_clk),
    .D(_01203_),
    .Q(\regs[27][19] ));
 sky130_fd_sc_hd__dfxtp_1 _15014_ (.CLK(clknet_leaf_13_clk),
    .D(_01204_),
    .Q(\regs[27][20] ));
 sky130_fd_sc_hd__dfxtp_1 _15015_ (.CLK(clknet_leaf_17_clk),
    .D(_01205_),
    .Q(\regs[27][21] ));
 sky130_fd_sc_hd__dfxtp_1 _15016_ (.CLK(clknet_leaf_117_clk),
    .D(_01206_),
    .Q(\regs[27][22] ));
 sky130_fd_sc_hd__dfxtp_1 _15017_ (.CLK(clknet_leaf_16_clk),
    .D(_01207_),
    .Q(\regs[27][23] ));
 sky130_fd_sc_hd__dfxtp_1 _15018_ (.CLK(clknet_leaf_15_clk),
    .D(_01208_),
    .Q(\regs[27][24] ));
 sky130_fd_sc_hd__dfxtp_1 _15019_ (.CLK(clknet_leaf_15_clk),
    .D(_01209_),
    .Q(\regs[27][25] ));
 sky130_fd_sc_hd__dfxtp_1 _15020_ (.CLK(clknet_leaf_18_clk),
    .D(_01210_),
    .Q(\regs[27][26] ));
 sky130_fd_sc_hd__dfxtp_1 _15021_ (.CLK(clknet_leaf_117_clk),
    .D(_01211_),
    .Q(\regs[27][27] ));
 sky130_fd_sc_hd__dfxtp_1 _15022_ (.CLK(clknet_leaf_12_clk),
    .D(_01212_),
    .Q(\regs[27][28] ));
 sky130_fd_sc_hd__dfxtp_1 _15023_ (.CLK(clknet_leaf_17_clk),
    .D(_01213_),
    .Q(\regs[27][29] ));
 sky130_fd_sc_hd__dfxtp_1 _15024_ (.CLK(clknet_leaf_116_clk),
    .D(_01214_),
    .Q(\regs[27][30] ));
 sky130_fd_sc_hd__dfxtp_1 _15025_ (.CLK(clknet_leaf_117_clk),
    .D(_01215_),
    .Q(\regs[27][31] ));
 sky130_fd_sc_hd__dfxtp_1 _15026_ (.CLK(clknet_leaf_15_clk),
    .D(_01216_),
    .Q(\regs[28][0] ));
 sky130_fd_sc_hd__dfxtp_1 _15027_ (.CLK(clknet_leaf_14_clk),
    .D(_01217_),
    .Q(\regs[28][1] ));
 sky130_fd_sc_hd__dfxtp_1 _15028_ (.CLK(clknet_leaf_121_clk),
    .D(_01218_),
    .Q(\regs[28][2] ));
 sky130_fd_sc_hd__dfxtp_1 _15029_ (.CLK(clknet_leaf_3_clk),
    .D(_01219_),
    .Q(\regs[28][3] ));
 sky130_fd_sc_hd__dfxtp_1 _15030_ (.CLK(clknet_leaf_119_clk),
    .D(_01220_),
    .Q(\regs[28][4] ));
 sky130_fd_sc_hd__dfxtp_1 _15031_ (.CLK(clknet_leaf_13_clk),
    .D(_01221_),
    .Q(\regs[28][5] ));
 sky130_fd_sc_hd__dfxtp_1 _15032_ (.CLK(clknet_leaf_108_clk),
    .D(_01222_),
    .Q(\regs[28][6] ));
 sky130_fd_sc_hd__dfxtp_1 _15033_ (.CLK(clknet_leaf_119_clk),
    .D(_01223_),
    .Q(\regs[28][7] ));
 sky130_fd_sc_hd__dfxtp_1 _15034_ (.CLK(clknet_leaf_3_clk),
    .D(_01224_),
    .Q(\regs[28][8] ));
 sky130_fd_sc_hd__dfxtp_1 _15035_ (.CLK(clknet_leaf_114_clk),
    .D(_01225_),
    .Q(\regs[28][9] ));
 sky130_fd_sc_hd__dfxtp_1 _15036_ (.CLK(clknet_leaf_111_clk),
    .D(_01226_),
    .Q(\regs[28][10] ));
 sky130_fd_sc_hd__dfxtp_1 _15037_ (.CLK(clknet_leaf_89_clk),
    .D(_01227_),
    .Q(\regs[28][11] ));
 sky130_fd_sc_hd__dfxtp_1 _15038_ (.CLK(clknet_leaf_88_clk),
    .D(_01228_),
    .Q(\regs[28][12] ));
 sky130_fd_sc_hd__dfxtp_1 _15039_ (.CLK(clknet_leaf_89_clk),
    .D(_01229_),
    .Q(\regs[28][13] ));
 sky130_fd_sc_hd__dfxtp_1 _15040_ (.CLK(clknet_leaf_82_clk),
    .D(_01230_),
    .Q(\regs[28][14] ));
 sky130_fd_sc_hd__dfxtp_1 _15041_ (.CLK(clknet_leaf_113_clk),
    .D(_01231_),
    .Q(\regs[28][15] ));
 sky130_fd_sc_hd__dfxtp_1 _15042_ (.CLK(clknet_leaf_89_clk),
    .D(_01232_),
    .Q(\regs[28][16] ));
 sky130_fd_sc_hd__dfxtp_1 _15043_ (.CLK(clknet_leaf_80_clk),
    .D(_01233_),
    .Q(\regs[28][17] ));
 sky130_fd_sc_hd__dfxtp_1 _15044_ (.CLK(clknet_leaf_112_clk),
    .D(_01234_),
    .Q(\regs[28][18] ));
 sky130_fd_sc_hd__dfxtp_1 _15045_ (.CLK(clknet_leaf_88_clk),
    .D(_01235_),
    .Q(\regs[28][19] ));
 sky130_fd_sc_hd__dfxtp_1 _15046_ (.CLK(clknet_leaf_11_clk),
    .D(_01236_),
    .Q(\regs[28][20] ));
 sky130_fd_sc_hd__dfxtp_1 _15047_ (.CLK(clknet_leaf_19_clk),
    .D(_01237_),
    .Q(\regs[28][21] ));
 sky130_fd_sc_hd__dfxtp_1 _15048_ (.CLK(clknet_leaf_19_clk),
    .D(_01238_),
    .Q(\regs[28][22] ));
 sky130_fd_sc_hd__dfxtp_1 _15049_ (.CLK(clknet_leaf_26_clk),
    .D(_01239_),
    .Q(\regs[28][23] ));
 sky130_fd_sc_hd__dfxtp_1 _15050_ (.CLK(clknet_leaf_21_clk),
    .D(_01240_),
    .Q(\regs[28][24] ));
 sky130_fd_sc_hd__dfxtp_1 _15051_ (.CLK(clknet_leaf_16_clk),
    .D(_01241_),
    .Q(\regs[28][25] ));
 sky130_fd_sc_hd__dfxtp_1 _15052_ (.CLK(clknet_leaf_19_clk),
    .D(_01242_),
    .Q(\regs[28][26] ));
 sky130_fd_sc_hd__dfxtp_1 _15053_ (.CLK(clknet_leaf_55_clk),
    .D(_01243_),
    .Q(\regs[28][27] ));
 sky130_fd_sc_hd__dfxtp_1 _15054_ (.CLK(clknet_leaf_11_clk),
    .D(_01244_),
    .Q(\regs[28][28] ));
 sky130_fd_sc_hd__dfxtp_1 _15055_ (.CLK(clknet_leaf_19_clk),
    .D(_01245_),
    .Q(\regs[28][29] ));
 sky130_fd_sc_hd__dfxtp_1 _15056_ (.CLK(clknet_leaf_116_clk),
    .D(_01246_),
    .Q(\regs[28][30] ));
 sky130_fd_sc_hd__dfxtp_1 _15057_ (.CLK(clknet_leaf_74_clk),
    .D(_01247_),
    .Q(\regs[28][31] ));
 sky130_fd_sc_hd__dfxtp_1 _15058_ (.CLK(clknet_leaf_131_clk),
    .D(_01248_),
    .Q(\regs[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _15059_ (.CLK(clknet_leaf_134_clk),
    .D(_01249_),
    .Q(\regs[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _15060_ (.CLK(clknet_leaf_129_clk),
    .D(_01250_),
    .Q(\regs[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _15061_ (.CLK(clknet_leaf_135_clk),
    .D(_01251_),
    .Q(\regs[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _15062_ (.CLK(clknet_leaf_130_clk),
    .D(_01252_),
    .Q(\regs[2][4] ));
 sky130_fd_sc_hd__dfxtp_1 _15063_ (.CLK(clknet_leaf_0_clk),
    .D(_01253_),
    .Q(\regs[2][5] ));
 sky130_fd_sc_hd__dfxtp_1 _15064_ (.CLK(clknet_leaf_126_clk),
    .D(_01254_),
    .Q(\regs[2][6] ));
 sky130_fd_sc_hd__dfxtp_1 _15065_ (.CLK(clknet_leaf_127_clk),
    .D(_01255_),
    .Q(\regs[2][7] ));
 sky130_fd_sc_hd__dfxtp_1 _15066_ (.CLK(clknet_leaf_0_clk),
    .D(_01256_),
    .Q(\regs[2][8] ));
 sky130_fd_sc_hd__dfxtp_1 _15067_ (.CLK(clknet_leaf_106_clk),
    .D(_01257_),
    .Q(\regs[2][9] ));
 sky130_fd_sc_hd__dfxtp_1 _15068_ (.CLK(clknet_leaf_101_clk),
    .D(_01258_),
    .Q(\regs[2][10] ));
 sky130_fd_sc_hd__dfxtp_1 _15069_ (.CLK(clknet_leaf_95_clk),
    .D(_01259_),
    .Q(\regs[2][11] ));
 sky130_fd_sc_hd__dfxtp_1 _15070_ (.CLK(clknet_leaf_101_clk),
    .D(_01260_),
    .Q(\regs[2][12] ));
 sky130_fd_sc_hd__dfxtp_1 _15071_ (.CLK(clknet_leaf_88_clk),
    .D(_01261_),
    .Q(\regs[2][13] ));
 sky130_fd_sc_hd__dfxtp_1 _15072_ (.CLK(clknet_leaf_94_clk),
    .D(_01262_),
    .Q(\regs[2][14] ));
 sky130_fd_sc_hd__dfxtp_1 _15073_ (.CLK(clknet_leaf_109_clk),
    .D(_01263_),
    .Q(\regs[2][15] ));
 sky130_fd_sc_hd__dfxtp_1 _15074_ (.CLK(clknet_leaf_94_clk),
    .D(_01264_),
    .Q(\regs[2][16] ));
 sky130_fd_sc_hd__dfxtp_1 _15075_ (.CLK(clknet_leaf_100_clk),
    .D(_01265_),
    .Q(\regs[2][17] ));
 sky130_fd_sc_hd__dfxtp_1 _15076_ (.CLK(clknet_leaf_110_clk),
    .D(_01266_),
    .Q(\regs[2][18] ));
 sky130_fd_sc_hd__dfxtp_1 _15077_ (.CLK(clknet_leaf_93_clk),
    .D(_01267_),
    .Q(\regs[2][19] ));
 sky130_fd_sc_hd__dfxtp_1 _15078_ (.CLK(clknet_leaf_8_clk),
    .D(_01268_),
    .Q(\regs[2][20] ));
 sky130_fd_sc_hd__dfxtp_1 _15079_ (.CLK(clknet_leaf_64_clk),
    .D(_01269_),
    .Q(\regs[2][21] ));
 sky130_fd_sc_hd__dfxtp_1 _15080_ (.CLK(clknet_leaf_64_clk),
    .D(_01270_),
    .Q(\regs[2][22] ));
 sky130_fd_sc_hd__dfxtp_1 _15081_ (.CLK(clknet_leaf_29_clk),
    .D(_01271_),
    .Q(\regs[2][23] ));
 sky130_fd_sc_hd__dfxtp_1 _15082_ (.CLK(clknet_leaf_26_clk),
    .D(_01272_),
    .Q(\regs[2][24] ));
 sky130_fd_sc_hd__dfxtp_1 _15083_ (.CLK(clknet_leaf_8_clk),
    .D(_01273_),
    .Q(\regs[2][25] ));
 sky130_fd_sc_hd__dfxtp_1 _15084_ (.CLK(clknet_leaf_69_clk),
    .D(_01274_),
    .Q(\regs[2][26] ));
 sky130_fd_sc_hd__dfxtp_1 _15085_ (.CLK(clknet_leaf_66_clk),
    .D(_01275_),
    .Q(\regs[2][27] ));
 sky130_fd_sc_hd__dfxtp_1 _15086_ (.CLK(clknet_leaf_29_clk),
    .D(_01276_),
    .Q(\regs[2][28] ));
 sky130_fd_sc_hd__dfxtp_1 _15087_ (.CLK(clknet_leaf_71_clk),
    .D(_01277_),
    .Q(\regs[2][29] ));
 sky130_fd_sc_hd__dfxtp_1 _15088_ (.CLK(clknet_leaf_73_clk),
    .D(_01278_),
    .Q(\regs[2][30] ));
 sky130_fd_sc_hd__dfxtp_1 _15089_ (.CLK(clknet_leaf_74_clk),
    .D(_01279_),
    .Q(\regs[2][31] ));
 sky130_fd_sc_hd__dfxtp_1 _15090_ (.CLK(clknet_leaf_15_clk),
    .D(_01280_),
    .Q(\regs[30][0] ));
 sky130_fd_sc_hd__dfxtp_1 _15091_ (.CLK(clknet_leaf_14_clk),
    .D(_01281_),
    .Q(\regs[30][1] ));
 sky130_fd_sc_hd__dfxtp_1 _15092_ (.CLK(clknet_leaf_121_clk),
    .D(_01282_),
    .Q(\regs[30][2] ));
 sky130_fd_sc_hd__dfxtp_1 _15093_ (.CLK(clknet_leaf_3_clk),
    .D(_01283_),
    .Q(\regs[30][3] ));
 sky130_fd_sc_hd__dfxtp_1 _15094_ (.CLK(clknet_leaf_121_clk),
    .D(_01284_),
    .Q(\regs[30][4] ));
 sky130_fd_sc_hd__dfxtp_1 _15095_ (.CLK(clknet_leaf_4_clk),
    .D(_01285_),
    .Q(\regs[30][5] ));
 sky130_fd_sc_hd__dfxtp_1 _15096_ (.CLK(clknet_leaf_108_clk),
    .D(_01286_),
    .Q(\regs[30][6] ));
 sky130_fd_sc_hd__dfxtp_1 _15097_ (.CLK(clknet_leaf_119_clk),
    .D(_01287_),
    .Q(\regs[30][7] ));
 sky130_fd_sc_hd__dfxtp_1 _15098_ (.CLK(clknet_leaf_3_clk),
    .D(_01288_),
    .Q(\regs[30][8] ));
 sky130_fd_sc_hd__dfxtp_1 _15099_ (.CLK(clknet_leaf_118_clk),
    .D(_01289_),
    .Q(\regs[30][9] ));
 sky130_fd_sc_hd__dfxtp_1 _15100_ (.CLK(clknet_leaf_111_clk),
    .D(_01290_),
    .Q(\regs[30][10] ));
 sky130_fd_sc_hd__dfxtp_1 _15101_ (.CLK(clknet_leaf_88_clk),
    .D(_01291_),
    .Q(\regs[30][11] ));
 sky130_fd_sc_hd__dfxtp_1 _15102_ (.CLK(clknet_leaf_90_clk),
    .D(_01292_),
    .Q(\regs[30][12] ));
 sky130_fd_sc_hd__dfxtp_1 _15103_ (.CLK(clknet_leaf_88_clk),
    .D(_01293_),
    .Q(\regs[30][13] ));
 sky130_fd_sc_hd__dfxtp_1 _15104_ (.CLK(clknet_leaf_83_clk),
    .D(_01294_),
    .Q(\regs[30][14] ));
 sky130_fd_sc_hd__dfxtp_1 _15105_ (.CLK(clknet_leaf_113_clk),
    .D(_01295_),
    .Q(\regs[30][15] ));
 sky130_fd_sc_hd__dfxtp_1 _15106_ (.CLK(clknet_leaf_88_clk),
    .D(_01296_),
    .Q(\regs[30][16] ));
 sky130_fd_sc_hd__dfxtp_1 _15107_ (.CLK(clknet_leaf_80_clk),
    .D(_01297_),
    .Q(\regs[30][17] ));
 sky130_fd_sc_hd__dfxtp_1 _15108_ (.CLK(clknet_leaf_78_clk),
    .D(_01298_),
    .Q(\regs[30][18] ));
 sky130_fd_sc_hd__dfxtp_1 _15109_ (.CLK(clknet_leaf_89_clk),
    .D(_01299_),
    .Q(\regs[30][19] ));
 sky130_fd_sc_hd__dfxtp_1 _15110_ (.CLK(clknet_leaf_10_clk),
    .D(_01300_),
    .Q(\regs[30][20] ));
 sky130_fd_sc_hd__dfxtp_1 _15111_ (.CLK(clknet_leaf_17_clk),
    .D(_01301_),
    .Q(\regs[30][21] ));
 sky130_fd_sc_hd__dfxtp_1 _15112_ (.CLK(clknet_leaf_19_clk),
    .D(_01302_),
    .Q(\regs[30][22] ));
 sky130_fd_sc_hd__dfxtp_1 _15113_ (.CLK(clknet_leaf_21_clk),
    .D(_01303_),
    .Q(\regs[30][23] ));
 sky130_fd_sc_hd__dfxtp_1 _15114_ (.CLK(clknet_leaf_21_clk),
    .D(_01304_),
    .Q(\regs[30][24] ));
 sky130_fd_sc_hd__dfxtp_1 _15115_ (.CLK(clknet_leaf_16_clk),
    .D(_01305_),
    .Q(\regs[30][25] ));
 sky130_fd_sc_hd__dfxtp_1 _15116_ (.CLK(clknet_leaf_19_clk),
    .D(_01306_),
    .Q(\regs[30][26] ));
 sky130_fd_sc_hd__dfxtp_1 _15117_ (.CLK(clknet_leaf_55_clk),
    .D(_01307_),
    .Q(\regs[30][27] ));
 sky130_fd_sc_hd__dfxtp_1 _15118_ (.CLK(clknet_leaf_10_clk),
    .D(_01308_),
    .Q(\regs[30][28] ));
 sky130_fd_sc_hd__dfxtp_1 _15119_ (.CLK(clknet_leaf_20_clk),
    .D(_01309_),
    .Q(\regs[30][29] ));
 sky130_fd_sc_hd__dfxtp_1 _15120_ (.CLK(clknet_leaf_115_clk),
    .D(_01310_),
    .Q(\regs[30][30] ));
 sky130_fd_sc_hd__dfxtp_1 _15121_ (.CLK(clknet_leaf_74_clk),
    .D(_01311_),
    .Q(\regs[30][31] ));
 sky130_fd_sc_hd__dfrtp_4 _15122_ (.CLK(clknet_leaf_124_clk),
    .D(_01312_),
    .RESET_B(_00073_),
    .Q(\rs2_content[0] ));
 sky130_fd_sc_hd__dfrtp_4 _15123_ (.CLK(clknet_leaf_118_clk),
    .D(_01313_),
    .RESET_B(_00074_),
    .Q(\rs2_content[1] ));
 sky130_fd_sc_hd__dfrtp_1 _15124_ (.CLK(clknet_leaf_53_clk),
    .D(_01314_),
    .RESET_B(_00075_),
    .Q(\rs2_content[2] ));
 sky130_fd_sc_hd__dfrtp_1 _15125_ (.CLK(clknet_leaf_57_clk),
    .D(_01315_),
    .RESET_B(_00076_),
    .Q(\rs2_content[3] ));
 sky130_fd_sc_hd__dfrtp_4 _15126_ (.CLK(clknet_leaf_123_clk),
    .D(_01316_),
    .RESET_B(_00077_),
    .Q(\rs2_content[4] ));
 sky130_fd_sc_hd__dfrtp_4 _15127_ (.CLK(clknet_leaf_118_clk),
    .D(_01317_),
    .RESET_B(_00078_),
    .Q(\rs2_content[5] ));
 sky130_fd_sc_hd__dfrtp_4 _15128_ (.CLK(clknet_leaf_109_clk),
    .D(_01318_),
    .RESET_B(_00079_),
    .Q(\rs2_content[6] ));
 sky130_fd_sc_hd__dfrtp_4 _15129_ (.CLK(clknet_leaf_108_clk),
    .D(_01319_),
    .RESET_B(_00080_),
    .Q(\rs2_content[7] ));
 sky130_fd_sc_hd__dfrtp_4 _15130_ (.CLK(clknet_leaf_114_clk),
    .D(_01320_),
    .RESET_B(_00081_),
    .Q(\rs2_content[8] ));
 sky130_fd_sc_hd__dfrtp_4 _15131_ (.CLK(clknet_leaf_109_clk),
    .D(_01321_),
    .RESET_B(_00082_),
    .Q(\rs2_content[9] ));
 sky130_fd_sc_hd__dfrtp_4 _15132_ (.CLK(clknet_leaf_78_clk),
    .D(_01322_),
    .RESET_B(_00083_),
    .Q(\rs2_content[10] ));
 sky130_fd_sc_hd__dfrtp_4 _15133_ (.CLK(clknet_leaf_89_clk),
    .D(_01323_),
    .RESET_B(_00084_),
    .Q(\rs2_content[11] ));
 sky130_fd_sc_hd__dfrtp_4 _15134_ (.CLK(clknet_leaf_90_clk),
    .D(_01324_),
    .RESET_B(_00085_),
    .Q(\rs2_content[12] ));
 sky130_fd_sc_hd__dfrtp_4 _15135_ (.CLK(clknet_leaf_79_clk),
    .D(_01325_),
    .RESET_B(_00086_),
    .Q(\rs2_content[13] ));
 sky130_fd_sc_hd__dfrtp_4 _15136_ (.CLK(clknet_leaf_82_clk),
    .D(_01326_),
    .RESET_B(_00087_),
    .Q(\rs2_content[14] ));
 sky130_fd_sc_hd__dfrtp_4 _15137_ (.CLK(clknet_leaf_76_clk),
    .D(_01327_),
    .RESET_B(_00088_),
    .Q(\rs2_content[15] ));
 sky130_fd_sc_hd__dfrtp_4 _15138_ (.CLK(clknet_leaf_82_clk),
    .D(_01328_),
    .RESET_B(_00089_),
    .Q(\rs2_content[16] ));
 sky130_fd_sc_hd__dfrtp_4 _15139_ (.CLK(clknet_leaf_81_clk),
    .D(_01329_),
    .RESET_B(_00090_),
    .Q(\rs2_content[17] ));
 sky130_fd_sc_hd__dfrtp_2 _15140_ (.CLK(clknet_leaf_81_clk),
    .D(_01330_),
    .RESET_B(_00091_),
    .Q(\rs2_content[18] ));
 sky130_fd_sc_hd__dfrtp_4 _15141_ (.CLK(clknet_leaf_82_clk),
    .D(_01331_),
    .RESET_B(_00092_),
    .Q(\rs2_content[19] ));
 sky130_fd_sc_hd__dfrtp_2 _15142_ (.CLK(clknet_leaf_67_clk),
    .D(_01332_),
    .RESET_B(_00093_),
    .Q(\rs2_content[20] ));
 sky130_fd_sc_hd__dfrtp_2 _15143_ (.CLK(clknet_leaf_64_clk),
    .D(_01333_),
    .RESET_B(_00094_),
    .Q(\rs2_content[21] ));
 sky130_fd_sc_hd__dfrtp_2 _15144_ (.CLK(clknet_leaf_64_clk),
    .D(_01334_),
    .RESET_B(_00095_),
    .Q(\rs2_content[22] ));
 sky130_fd_sc_hd__dfrtp_1 _15145_ (.CLK(clknet_leaf_67_clk),
    .D(_01335_),
    .RESET_B(_00096_),
    .Q(\rs2_content[23] ));
 sky130_fd_sc_hd__dfrtp_4 _15146_ (.CLK(clknet_leaf_56_clk),
    .D(_01336_),
    .RESET_B(_00097_),
    .Q(\rs2_content[24] ));
 sky130_fd_sc_hd__dfrtp_2 _15147_ (.CLK(clknet_leaf_62_clk),
    .D(_01337_),
    .RESET_B(_00098_),
    .Q(\rs2_content[25] ));
 sky130_fd_sc_hd__dfrtp_1 _15148_ (.CLK(clknet_leaf_68_clk),
    .D(_01338_),
    .RESET_B(_00099_),
    .Q(\rs2_content[26] ));
 sky130_fd_sc_hd__dfrtp_2 _15149_ (.CLK(clknet_leaf_68_clk),
    .D(_01339_),
    .RESET_B(_00100_),
    .Q(\rs2_content[27] ));
 sky130_fd_sc_hd__dfrtp_4 _15150_ (.CLK(clknet_leaf_25_clk),
    .D(_01340_),
    .RESET_B(_00101_),
    .Q(\rs2_content[28] ));
 sky130_fd_sc_hd__dfrtp_2 _15151_ (.CLK(clknet_leaf_68_clk),
    .D(_01341_),
    .RESET_B(_00102_),
    .Q(\rs2_content[29] ));
 sky130_fd_sc_hd__dfrtp_4 _15152_ (.CLK(clknet_leaf_56_clk),
    .D(_01342_),
    .RESET_B(_00103_),
    .Q(\rs2_content[30] ));
 sky130_fd_sc_hd__dfrtp_2 _15153_ (.CLK(clknet_leaf_68_clk),
    .D(_01343_),
    .RESET_B(_00104_),
    .Q(\rs2_content[31] ));
 sky130_fd_sc_hd__dfrtp_1 _15154_ (.CLK(clknet_leaf_25_clk),
    .D(_01344_),
    .RESET_B(_00105_),
    .Q(\instret[0] ));
 sky130_fd_sc_hd__dfrtp_1 _15155_ (.CLK(clknet_leaf_25_clk),
    .D(_01345_),
    .RESET_B(_00106_),
    .Q(\instret[1] ));
 sky130_fd_sc_hd__dfrtp_1 _15156_ (.CLK(clknet_leaf_25_clk),
    .D(_01346_),
    .RESET_B(_00107_),
    .Q(\instret[2] ));
 sky130_fd_sc_hd__dfrtp_1 _15157_ (.CLK(clknet_leaf_24_clk),
    .D(_01347_),
    .RESET_B(_00108_),
    .Q(\instret[3] ));
 sky130_fd_sc_hd__dfrtp_1 _15158_ (.CLK(clknet_leaf_33_clk),
    .D(_01348_),
    .RESET_B(_00109_),
    .Q(\instret[4] ));
 sky130_fd_sc_hd__dfrtp_1 _15159_ (.CLK(clknet_leaf_33_clk),
    .D(_01349_),
    .RESET_B(_00110_),
    .Q(\instret[5] ));
 sky130_fd_sc_hd__dfrtp_1 _15160_ (.CLK(clknet_leaf_33_clk),
    .D(_01350_),
    .RESET_B(_00111_),
    .Q(\instret[6] ));
 sky130_fd_sc_hd__dfrtp_1 _15161_ (.CLK(clknet_leaf_33_clk),
    .D(_01351_),
    .RESET_B(_00112_),
    .Q(\instret[7] ));
 sky130_fd_sc_hd__dfrtp_1 _15162_ (.CLK(clknet_leaf_33_clk),
    .D(_01352_),
    .RESET_B(_00113_),
    .Q(\instret[8] ));
 sky130_fd_sc_hd__dfrtp_1 _15163_ (.CLK(clknet_leaf_33_clk),
    .D(_01353_),
    .RESET_B(_00114_),
    .Q(\instret[9] ));
 sky130_fd_sc_hd__dfrtp_1 _15164_ (.CLK(clknet_leaf_34_clk),
    .D(_01354_),
    .RESET_B(_00115_),
    .Q(\instret[10] ));
 sky130_fd_sc_hd__dfrtp_1 _15165_ (.CLK(clknet_leaf_41_clk),
    .D(_01355_),
    .RESET_B(_00116_),
    .Q(\instret[11] ));
 sky130_fd_sc_hd__dfrtp_1 _15166_ (.CLK(clknet_leaf_41_clk),
    .D(_01356_),
    .RESET_B(_00117_),
    .Q(\instret[12] ));
 sky130_fd_sc_hd__dfrtp_1 _15167_ (.CLK(clknet_leaf_41_clk),
    .D(_01357_),
    .RESET_B(_00118_),
    .Q(\instret[13] ));
 sky130_fd_sc_hd__dfrtp_1 _15168_ (.CLK(clknet_leaf_41_clk),
    .D(_01358_),
    .RESET_B(_00119_),
    .Q(\instret[14] ));
 sky130_fd_sc_hd__dfrtp_1 _15169_ (.CLK(clknet_leaf_41_clk),
    .D(_01359_),
    .RESET_B(_00120_),
    .Q(\instret[15] ));
 sky130_fd_sc_hd__dfrtp_1 _15170_ (.CLK(clknet_leaf_40_clk),
    .D(_01360_),
    .RESET_B(_00121_),
    .Q(\instret[16] ));
 sky130_fd_sc_hd__dfrtp_1 _15171_ (.CLK(clknet_leaf_40_clk),
    .D(_01361_),
    .RESET_B(_00122_),
    .Q(\instret[17] ));
 sky130_fd_sc_hd__dfrtp_1 _15172_ (.CLK(clknet_leaf_40_clk),
    .D(_01362_),
    .RESET_B(_00123_),
    .Q(\instret[18] ));
 sky130_fd_sc_hd__dfrtp_1 _15173_ (.CLK(clknet_leaf_43_clk),
    .D(_01363_),
    .RESET_B(_00124_),
    .Q(\instret[19] ));
 sky130_fd_sc_hd__dfrtp_1 _15174_ (.CLK(clknet_leaf_43_clk),
    .D(_01364_),
    .RESET_B(_00125_),
    .Q(\instret[20] ));
 sky130_fd_sc_hd__dfrtp_1 _15175_ (.CLK(clknet_leaf_43_clk),
    .D(_01365_),
    .RESET_B(_00126_),
    .Q(\instret[21] ));
 sky130_fd_sc_hd__dfrtp_1 _15176_ (.CLK(clknet_leaf_40_clk),
    .D(_01366_),
    .RESET_B(_00127_),
    .Q(\instret[22] ));
 sky130_fd_sc_hd__dfrtp_1 _15177_ (.CLK(clknet_leaf_41_clk),
    .D(_01367_),
    .RESET_B(_00128_),
    .Q(\instret[23] ));
 sky130_fd_sc_hd__dfrtp_1 _15178_ (.CLK(clknet_leaf_42_clk),
    .D(_01368_),
    .RESET_B(_00129_),
    .Q(\instret[24] ));
 sky130_fd_sc_hd__dfrtp_1 _15179_ (.CLK(clknet_leaf_42_clk),
    .D(_01369_),
    .RESET_B(_00130_),
    .Q(\instret[25] ));
 sky130_fd_sc_hd__dfrtp_1 _15180_ (.CLK(clknet_leaf_42_clk),
    .D(_01370_),
    .RESET_B(_00131_),
    .Q(\instret[26] ));
 sky130_fd_sc_hd__dfrtp_1 _15181_ (.CLK(clknet_leaf_33_clk),
    .D(_01371_),
    .RESET_B(_00132_),
    .Q(\instret[27] ));
 sky130_fd_sc_hd__dfrtp_1 _15182_ (.CLK(clknet_leaf_33_clk),
    .D(_01372_),
    .RESET_B(_00133_),
    .Q(\instret[28] ));
 sky130_fd_sc_hd__dfrtp_1 _15183_ (.CLK(clknet_leaf_33_clk),
    .D(_01373_),
    .RESET_B(_00134_),
    .Q(\instret[29] ));
 sky130_fd_sc_hd__dfrtp_1 _15184_ (.CLK(clknet_leaf_24_clk),
    .D(_01374_),
    .RESET_B(_00135_),
    .Q(\instret[30] ));
 sky130_fd_sc_hd__dfrtp_1 _15185_ (.CLK(clknet_leaf_24_clk),
    .D(_01375_),
    .RESET_B(_00136_),
    .Q(\instret[31] ));
 sky130_fd_sc_hd__dfrtp_1 _15186_ (.CLK(clknet_leaf_24_clk),
    .D(_01376_),
    .RESET_B(_00137_),
    .Q(\instret[32] ));
 sky130_fd_sc_hd__dfrtp_1 _15187_ (.CLK(clknet_leaf_32_clk),
    .D(_01377_),
    .RESET_B(_00138_),
    .Q(\instret[33] ));
 sky130_fd_sc_hd__dfrtp_1 _15188_ (.CLK(clknet_leaf_32_clk),
    .D(_01378_),
    .RESET_B(_00139_),
    .Q(\instret[34] ));
 sky130_fd_sc_hd__dfrtp_1 _15189_ (.CLK(clknet_leaf_32_clk),
    .D(_01379_),
    .RESET_B(_00140_),
    .Q(\instret[35] ));
 sky130_fd_sc_hd__dfrtp_1 _15190_ (.CLK(clknet_leaf_32_clk),
    .D(_01380_),
    .RESET_B(_00141_),
    .Q(\instret[36] ));
 sky130_fd_sc_hd__dfrtp_1 _15191_ (.CLK(clknet_leaf_32_clk),
    .D(_01381_),
    .RESET_B(_00142_),
    .Q(\instret[37] ));
 sky130_fd_sc_hd__dfrtp_1 _15192_ (.CLK(clknet_leaf_33_clk),
    .D(_01382_),
    .RESET_B(_00143_),
    .Q(\instret[38] ));
 sky130_fd_sc_hd__dfrtp_1 _15193_ (.CLK(clknet_leaf_33_clk),
    .D(_01383_),
    .RESET_B(_00144_),
    .Q(\instret[39] ));
 sky130_fd_sc_hd__dfrtp_1 _15194_ (.CLK(clknet_leaf_34_clk),
    .D(_01384_),
    .RESET_B(_00145_),
    .Q(\instret[40] ));
 sky130_fd_sc_hd__dfrtp_1 _15195_ (.CLK(clknet_leaf_34_clk),
    .D(_01385_),
    .RESET_B(_00146_),
    .Q(\instret[41] ));
 sky130_fd_sc_hd__dfrtp_1 _15196_ (.CLK(clknet_leaf_41_clk),
    .D(_01386_),
    .RESET_B(_00147_),
    .Q(\instret[42] ));
 sky130_fd_sc_hd__dfrtp_1 _15197_ (.CLK(clknet_leaf_41_clk),
    .D(_01387_),
    .RESET_B(_00148_),
    .Q(\instret[43] ));
 sky130_fd_sc_hd__dfrtp_1 _15198_ (.CLK(clknet_leaf_39_clk),
    .D(_01388_),
    .RESET_B(_00149_),
    .Q(\instret[44] ));
 sky130_fd_sc_hd__dfrtp_1 _15199_ (.CLK(clknet_leaf_39_clk),
    .D(_01389_),
    .RESET_B(_00150_),
    .Q(\instret[45] ));
 sky130_fd_sc_hd__dfrtp_1 _15200_ (.CLK(clknet_leaf_39_clk),
    .D(_01390_),
    .RESET_B(_00151_),
    .Q(\instret[46] ));
 sky130_fd_sc_hd__dfrtp_1 _15201_ (.CLK(clknet_leaf_39_clk),
    .D(_01391_),
    .RESET_B(_00152_),
    .Q(\instret[47] ));
 sky130_fd_sc_hd__dfrtp_1 _15202_ (.CLK(clknet_leaf_39_clk),
    .D(_01392_),
    .RESET_B(_00153_),
    .Q(\instret[48] ));
 sky130_fd_sc_hd__dfrtp_1 _15203_ (.CLK(clknet_leaf_39_clk),
    .D(_01393_),
    .RESET_B(_00154_),
    .Q(\instret[49] ));
 sky130_fd_sc_hd__dfrtp_1 _15204_ (.CLK(clknet_leaf_39_clk),
    .D(_01394_),
    .RESET_B(_00155_),
    .Q(\instret[50] ));
 sky130_fd_sc_hd__dfrtp_1 _15205_ (.CLK(clknet_leaf_39_clk),
    .D(_01395_),
    .RESET_B(_00156_),
    .Q(\instret[51] ));
 sky130_fd_sc_hd__dfrtp_1 _15206_ (.CLK(clknet_leaf_40_clk),
    .D(_01396_),
    .RESET_B(_00157_),
    .Q(\instret[52] ));
 sky130_fd_sc_hd__dfrtp_1 _15207_ (.CLK(clknet_leaf_44_clk),
    .D(_01397_),
    .RESET_B(_00158_),
    .Q(\instret[53] ));
 sky130_fd_sc_hd__dfrtp_1 _15208_ (.CLK(clknet_leaf_42_clk),
    .D(_01398_),
    .RESET_B(_00159_),
    .Q(\instret[54] ));
 sky130_fd_sc_hd__dfrtp_1 _15209_ (.CLK(clknet_leaf_42_clk),
    .D(_01399_),
    .RESET_B(_00160_),
    .Q(\instret[55] ));
 sky130_fd_sc_hd__dfrtp_1 _15210_ (.CLK(clknet_leaf_42_clk),
    .D(_01400_),
    .RESET_B(_00161_),
    .Q(\instret[56] ));
 sky130_fd_sc_hd__dfrtp_1 _15211_ (.CLK(clknet_leaf_42_clk),
    .D(_01401_),
    .RESET_B(_00162_),
    .Q(\instret[57] ));
 sky130_fd_sc_hd__dfrtp_1 _15212_ (.CLK(clknet_leaf_42_clk),
    .D(_01402_),
    .RESET_B(_00163_),
    .Q(\instret[58] ));
 sky130_fd_sc_hd__dfrtp_1 _15213_ (.CLK(clknet_leaf_42_clk),
    .D(_01403_),
    .RESET_B(_00164_),
    .Q(\instret[59] ));
 sky130_fd_sc_hd__dfrtp_1 _15214_ (.CLK(clknet_leaf_42_clk),
    .D(_01404_),
    .RESET_B(_00165_),
    .Q(\instret[60] ));
 sky130_fd_sc_hd__dfrtp_1 _15215_ (.CLK(clknet_leaf_50_clk),
    .D(_01405_),
    .RESET_B(_00166_),
    .Q(\instret[61] ));
 sky130_fd_sc_hd__dfrtp_1 _15216_ (.CLK(clknet_leaf_50_clk),
    .D(_01406_),
    .RESET_B(_00167_),
    .Q(\instret[62] ));
 sky130_fd_sc_hd__dfrtp_1 _15217_ (.CLK(clknet_leaf_50_clk),
    .D(_01407_),
    .RESET_B(_00168_),
    .Q(\instret[63] ));
 sky130_fd_sc_hd__dfrtp_4 _15218_ (.CLK(clknet_leaf_52_clk),
    .D(_01408_),
    .RESET_B(_00169_),
    .Q(\leorv32_alu.input1[0] ));
 sky130_fd_sc_hd__dfrtp_4 _15219_ (.CLK(clknet_leaf_51_clk),
    .D(_01409_),
    .RESET_B(_00170_),
    .Q(\leorv32_alu.input1[1] ));
 sky130_fd_sc_hd__dfrtp_2 _15220_ (.CLK(clknet_leaf_57_clk),
    .D(_01410_),
    .RESET_B(_00171_),
    .Q(\leorv32_alu.input1[2] ));
 sky130_fd_sc_hd__dfrtp_1 _15221_ (.CLK(clknet_leaf_57_clk),
    .D(_01411_),
    .RESET_B(_00172_),
    .Q(\leorv32_alu.input1[3] ));
 sky130_fd_sc_hd__dfrtp_1 _15222_ (.CLK(clknet_leaf_52_clk),
    .D(_01412_),
    .RESET_B(_00173_),
    .Q(\leorv32_alu.input1[4] ));
 sky130_fd_sc_hd__dfrtp_4 _15223_ (.CLK(clknet_leaf_24_clk),
    .D(_01413_),
    .RESET_B(_00174_),
    .Q(\leorv32_alu.input1[5] ));
 sky130_fd_sc_hd__dfrtp_4 _15224_ (.CLK(clknet_leaf_56_clk),
    .D(_01414_),
    .RESET_B(_00175_),
    .Q(\leorv32_alu.input1[6] ));
 sky130_fd_sc_hd__dfrtp_1 _15225_ (.CLK(clknet_leaf_57_clk),
    .D(_01415_),
    .RESET_B(_00176_),
    .Q(\leorv32_alu.input1[7] ));
 sky130_fd_sc_hd__dfrtp_4 _15226_ (.CLK(clknet_leaf_24_clk),
    .D(_01416_),
    .RESET_B(_00177_),
    .Q(\leorv32_alu.input1[8] ));
 sky130_fd_sc_hd__dfrtp_1 _15227_ (.CLK(clknet_leaf_56_clk),
    .D(_01417_),
    .RESET_B(_00178_),
    .Q(\leorv32_alu.input1[9] ));
 sky130_fd_sc_hd__dfrtp_1 _15228_ (.CLK(clknet_leaf_68_clk),
    .D(_01418_),
    .RESET_B(_00179_),
    .Q(\leorv32_alu.input1[10] ));
 sky130_fd_sc_hd__dfrtp_1 _15229_ (.CLK(clknet_leaf_67_clk),
    .D(_01419_),
    .RESET_B(_00180_),
    .Q(\leorv32_alu.input1[11] ));
 sky130_fd_sc_hd__dfrtp_1 _15230_ (.CLK(clknet_leaf_67_clk),
    .D(_01420_),
    .RESET_B(_00181_),
    .Q(\leorv32_alu.input1[12] ));
 sky130_fd_sc_hd__dfrtp_1 _15231_ (.CLK(clknet_leaf_67_clk),
    .D(_01421_),
    .RESET_B(_00182_),
    .Q(\leorv32_alu.input1[13] ));
 sky130_fd_sc_hd__dfrtp_1 _15232_ (.CLK(clknet_leaf_67_clk),
    .D(_01422_),
    .RESET_B(_00183_),
    .Q(\leorv32_alu.input1[14] ));
 sky130_fd_sc_hd__dfrtp_2 _15233_ (.CLK(clknet_leaf_68_clk),
    .D(_01423_),
    .RESET_B(_00184_),
    .Q(\leorv32_alu.input1[15] ));
 sky130_fd_sc_hd__dfrtp_1 _15234_ (.CLK(clknet_leaf_67_clk),
    .D(_01424_),
    .RESET_B(_00185_),
    .Q(\leorv32_alu.input1[16] ));
 sky130_fd_sc_hd__dfrtp_1 _15235_ (.CLK(clknet_leaf_67_clk),
    .D(_01425_),
    .RESET_B(_00186_),
    .Q(\leorv32_alu.input1[17] ));
 sky130_fd_sc_hd__dfrtp_1 _15236_ (.CLK(clknet_leaf_67_clk),
    .D(_01426_),
    .RESET_B(_00187_),
    .Q(\leorv32_alu.input1[18] ));
 sky130_fd_sc_hd__dfrtp_1 _15237_ (.CLK(clknet_leaf_67_clk),
    .D(_01427_),
    .RESET_B(_00188_),
    .Q(\leorv32_alu.input1[19] ));
 sky130_fd_sc_hd__dfrtp_4 _15238_ (.CLK(clknet_leaf_56_clk),
    .D(_01428_),
    .RESET_B(_00189_),
    .Q(\leorv32_alu.input1[20] ));
 sky130_fd_sc_hd__dfrtp_4 _15239_ (.CLK(clknet_leaf_66_clk),
    .D(_01429_),
    .RESET_B(_00190_),
    .Q(\leorv32_alu.input1[21] ));
 sky130_fd_sc_hd__dfrtp_4 _15240_ (.CLK(clknet_leaf_66_clk),
    .D(_01430_),
    .RESET_B(_00191_),
    .Q(\leorv32_alu.input1[22] ));
 sky130_fd_sc_hd__dfrtp_4 _15241_ (.CLK(clknet_leaf_56_clk),
    .D(_01431_),
    .RESET_B(_00192_),
    .Q(\leorv32_alu.input1[23] ));
 sky130_fd_sc_hd__dfrtp_4 _15242_ (.CLK(clknet_leaf_56_clk),
    .D(_01432_),
    .RESET_B(_00193_),
    .Q(\leorv32_alu.input1[24] ));
 sky130_fd_sc_hd__dfrtp_4 _15243_ (.CLK(clknet_leaf_56_clk),
    .D(_01433_),
    .RESET_B(_00194_),
    .Q(\leorv32_alu.input1[25] ));
 sky130_fd_sc_hd__dfrtp_4 _15244_ (.CLK(clknet_leaf_69_clk),
    .D(_01434_),
    .RESET_B(_00195_),
    .Q(\leorv32_alu.input1[26] ));
 sky130_fd_sc_hd__dfrtp_4 _15245_ (.CLK(clknet_leaf_66_clk),
    .D(_01435_),
    .RESET_B(_00196_),
    .Q(\leorv32_alu.input1[27] ));
 sky130_fd_sc_hd__dfrtp_1 _15246_ (.CLK(clknet_leaf_68_clk),
    .D(_01436_),
    .RESET_B(_00197_),
    .Q(\leorv32_alu.input1[28] ));
 sky130_fd_sc_hd__dfrtp_4 _15247_ (.CLK(clknet_leaf_68_clk),
    .D(_01437_),
    .RESET_B(_00198_),
    .Q(\leorv32_alu.input1[29] ));
 sky130_fd_sc_hd__dfrtp_4 _15248_ (.CLK(clknet_leaf_56_clk),
    .D(_01438_),
    .RESET_B(_00199_),
    .Q(\leorv32_alu.input1[30] ));
 sky130_fd_sc_hd__dfrtp_4 _15249_ (.CLK(clknet_4_12_0_clk),
    .D(_01439_),
    .RESET_B(_00200_),
    .Q(\leorv32_alu.input1[31] ));
 sky130_fd_sc_hd__dfrtp_2 _15250_ (.CLK(clknet_leaf_25_clk),
    .D(_00004_),
    .RESET_B(_00201_),
    .Q(\cycles[0] ));
 sky130_fd_sc_hd__dfrtp_1 _15251_ (.CLK(clknet_leaf_25_clk),
    .D(_00015_),
    .RESET_B(_00202_),
    .Q(\cycles[1] ));
 sky130_fd_sc_hd__dfrtp_1 _15252_ (.CLK(clknet_leaf_32_clk),
    .D(_00026_),
    .RESET_B(_00203_),
    .Q(\cycles[2] ));
 sky130_fd_sc_hd__dfrtp_1 _15253_ (.CLK(clknet_leaf_32_clk),
    .D(_00037_),
    .RESET_B(_00204_),
    .Q(\cycles[3] ));
 sky130_fd_sc_hd__dfrtp_1 _15254_ (.CLK(clknet_leaf_32_clk),
    .D(_00048_),
    .RESET_B(_00205_),
    .Q(\cycles[4] ));
 sky130_fd_sc_hd__dfrtp_1 _15255_ (.CLK(clknet_leaf_32_clk),
    .D(_00059_),
    .RESET_B(_00206_),
    .Q(\cycles[5] ));
 sky130_fd_sc_hd__dfrtp_1 _15256_ (.CLK(clknet_leaf_32_clk),
    .D(_00064_),
    .RESET_B(_00207_),
    .Q(\cycles[6] ));
 sky130_fd_sc_hd__dfrtp_1 _15257_ (.CLK(clknet_leaf_34_clk),
    .D(_00065_),
    .RESET_B(_00208_),
    .Q(\cycles[7] ));
 sky130_fd_sc_hd__dfrtp_1 _15258_ (.CLK(clknet_leaf_34_clk),
    .D(_00066_),
    .RESET_B(_00209_),
    .Q(\cycles[8] ));
 sky130_fd_sc_hd__dfrtp_1 _15259_ (.CLK(clknet_leaf_34_clk),
    .D(_00067_),
    .RESET_B(_00210_),
    .Q(\cycles[9] ));
 sky130_fd_sc_hd__dfrtp_1 _15260_ (.CLK(clknet_leaf_34_clk),
    .D(_00005_),
    .RESET_B(_00211_),
    .Q(\cycles[10] ));
 sky130_fd_sc_hd__dfrtp_1 _15261_ (.CLK(clknet_leaf_34_clk),
    .D(_00006_),
    .RESET_B(_00212_),
    .Q(\cycles[11] ));
 sky130_fd_sc_hd__dfrtp_1 _15262_ (.CLK(clknet_leaf_34_clk),
    .D(_00007_),
    .RESET_B(_00213_),
    .Q(\cycles[12] ));
 sky130_fd_sc_hd__dfrtp_1 _15263_ (.CLK(clknet_leaf_34_clk),
    .D(_00008_),
    .RESET_B(_00214_),
    .Q(\cycles[13] ));
 sky130_fd_sc_hd__dfrtp_1 _15264_ (.CLK(clknet_leaf_41_clk),
    .D(_00009_),
    .RESET_B(_00215_),
    .Q(\cycles[14] ));
 sky130_fd_sc_hd__dfrtp_1 _15265_ (.CLK(clknet_leaf_37_clk),
    .D(_00010_),
    .RESET_B(_00216_),
    .Q(\cycles[15] ));
 sky130_fd_sc_hd__dfrtp_1 _15266_ (.CLK(clknet_leaf_38_clk),
    .D(_00011_),
    .RESET_B(_00217_),
    .Q(\cycles[16] ));
 sky130_fd_sc_hd__dfrtp_1 _15267_ (.CLK(clknet_leaf_38_clk),
    .D(_00012_),
    .RESET_B(_00218_),
    .Q(\cycles[17] ));
 sky130_fd_sc_hd__dfrtp_1 _15268_ (.CLK(clknet_leaf_37_clk),
    .D(_00013_),
    .RESET_B(_00219_),
    .Q(\cycles[18] ));
 sky130_fd_sc_hd__dfrtp_1 _15269_ (.CLK(clknet_leaf_37_clk),
    .D(_00014_),
    .RESET_B(_00220_),
    .Q(\cycles[19] ));
 sky130_fd_sc_hd__dfrtp_1 _15270_ (.CLK(clknet_leaf_37_clk),
    .D(_00016_),
    .RESET_B(_00221_),
    .Q(\cycles[20] ));
 sky130_fd_sc_hd__dfrtp_1 _15271_ (.CLK(clknet_leaf_37_clk),
    .D(_00017_),
    .RESET_B(_00222_),
    .Q(\cycles[21] ));
 sky130_fd_sc_hd__dfrtp_1 _15272_ (.CLK(clknet_leaf_36_clk),
    .D(_00018_),
    .RESET_B(_00223_),
    .Q(\cycles[22] ));
 sky130_fd_sc_hd__dfrtp_1 _15273_ (.CLK(clknet_leaf_36_clk),
    .D(_00019_),
    .RESET_B(_00224_),
    .Q(\cycles[23] ));
 sky130_fd_sc_hd__dfrtp_1 _15274_ (.CLK(clknet_leaf_36_clk),
    .D(_00020_),
    .RESET_B(_00225_),
    .Q(\cycles[24] ));
 sky130_fd_sc_hd__dfrtp_1 _15275_ (.CLK(clknet_leaf_35_clk),
    .D(_00021_),
    .RESET_B(_00226_),
    .Q(\cycles[25] ));
 sky130_fd_sc_hd__dfrtp_1 _15276_ (.CLK(clknet_leaf_35_clk),
    .D(_00022_),
    .RESET_B(_00227_),
    .Q(\cycles[26] ));
 sky130_fd_sc_hd__dfrtp_1 _15277_ (.CLK(clknet_leaf_35_clk),
    .D(_00023_),
    .RESET_B(_00228_),
    .Q(\cycles[27] ));
 sky130_fd_sc_hd__dfrtp_1 _15278_ (.CLK(clknet_leaf_35_clk),
    .D(_00024_),
    .RESET_B(_00229_),
    .Q(\cycles[28] ));
 sky130_fd_sc_hd__dfrtp_1 _15279_ (.CLK(clknet_leaf_31_clk),
    .D(_00025_),
    .RESET_B(_00230_),
    .Q(\cycles[29] ));
 sky130_fd_sc_hd__dfrtp_1 _15280_ (.CLK(clknet_leaf_31_clk),
    .D(_00027_),
    .RESET_B(_00231_),
    .Q(\cycles[30] ));
 sky130_fd_sc_hd__dfrtp_1 _15281_ (.CLK(clknet_leaf_31_clk),
    .D(_00028_),
    .RESET_B(_00232_),
    .Q(\cycles[31] ));
 sky130_fd_sc_hd__dfrtp_1 _15282_ (.CLK(clknet_leaf_31_clk),
    .D(_00029_),
    .RESET_B(_00233_),
    .Q(\cycles[32] ));
 sky130_fd_sc_hd__dfrtp_1 _15283_ (.CLK(clknet_leaf_32_clk),
    .D(_00030_),
    .RESET_B(_00234_),
    .Q(\cycles[33] ));
 sky130_fd_sc_hd__dfrtp_1 _15284_ (.CLK(clknet_leaf_32_clk),
    .D(_00031_),
    .RESET_B(_00235_),
    .Q(\cycles[34] ));
 sky130_fd_sc_hd__dfrtp_2 _15285_ (.CLK(clknet_leaf_31_clk),
    .D(_00032_),
    .RESET_B(_00236_),
    .Q(\cycles[35] ));
 sky130_fd_sc_hd__dfrtp_1 _15286_ (.CLK(clknet_leaf_31_clk),
    .D(_00033_),
    .RESET_B(_00237_),
    .Q(\cycles[36] ));
 sky130_fd_sc_hd__dfrtp_1 _15287_ (.CLK(clknet_leaf_31_clk),
    .D(_00034_),
    .RESET_B(_00238_),
    .Q(\cycles[37] ));
 sky130_fd_sc_hd__dfrtp_1 _15288_ (.CLK(clknet_leaf_31_clk),
    .D(_00035_),
    .RESET_B(_00239_),
    .Q(\cycles[38] ));
 sky130_fd_sc_hd__dfrtp_1 _15289_ (.CLK(clknet_leaf_35_clk),
    .D(_00036_),
    .RESET_B(_00240_),
    .Q(\cycles[39] ));
 sky130_fd_sc_hd__dfrtp_1 _15290_ (.CLK(clknet_leaf_35_clk),
    .D(_00038_),
    .RESET_B(_00241_),
    .Q(\cycles[40] ));
 sky130_fd_sc_hd__dfrtp_1 _15291_ (.CLK(clknet_leaf_35_clk),
    .D(_00039_),
    .RESET_B(_00242_),
    .Q(\cycles[41] ));
 sky130_fd_sc_hd__dfrtp_1 _15292_ (.CLK(clknet_leaf_34_clk),
    .D(_00040_),
    .RESET_B(_00243_),
    .Q(\cycles[42] ));
 sky130_fd_sc_hd__dfrtp_1 _15293_ (.CLK(clknet_leaf_34_clk),
    .D(_00041_),
    .RESET_B(_00244_),
    .Q(\cycles[43] ));
 sky130_fd_sc_hd__dfrtp_1 _15294_ (.CLK(clknet_leaf_36_clk),
    .D(_00042_),
    .RESET_B(_00245_),
    .Q(\cycles[44] ));
 sky130_fd_sc_hd__dfrtp_1 _15295_ (.CLK(clknet_leaf_36_clk),
    .D(_00043_),
    .RESET_B(_00246_),
    .Q(\cycles[45] ));
 sky130_fd_sc_hd__dfrtp_1 _15296_ (.CLK(clknet_leaf_36_clk),
    .D(_00044_),
    .RESET_B(_00247_),
    .Q(\cycles[46] ));
 sky130_fd_sc_hd__dfrtp_1 _15297_ (.CLK(clknet_leaf_37_clk),
    .D(_00045_),
    .RESET_B(_00248_),
    .Q(\cycles[47] ));
 sky130_fd_sc_hd__dfrtp_1 _15298_ (.CLK(clknet_leaf_38_clk),
    .D(_00046_),
    .RESET_B(_00249_),
    .Q(\cycles[48] ));
 sky130_fd_sc_hd__dfrtp_1 _15299_ (.CLK(clknet_leaf_38_clk),
    .D(_00047_),
    .RESET_B(_00250_),
    .Q(\cycles[49] ));
 sky130_fd_sc_hd__dfrtp_1 _15300_ (.CLK(clknet_leaf_37_clk),
    .D(_00049_),
    .RESET_B(_00251_),
    .Q(\cycles[50] ));
 sky130_fd_sc_hd__dfrtp_1 _15301_ (.CLK(clknet_leaf_37_clk),
    .D(_00050_),
    .RESET_B(_00252_),
    .Q(\cycles[51] ));
 sky130_fd_sc_hd__dfrtp_1 _15302_ (.CLK(clknet_leaf_38_clk),
    .D(_00051_),
    .RESET_B(_00253_),
    .Q(\cycles[52] ));
 sky130_fd_sc_hd__dfrtp_1 _15303_ (.CLK(clknet_leaf_38_clk),
    .D(_00052_),
    .RESET_B(_00254_),
    .Q(\cycles[53] ));
 sky130_fd_sc_hd__dfrtp_1 _15304_ (.CLK(clknet_leaf_36_clk),
    .D(_00053_),
    .RESET_B(_00255_),
    .Q(\cycles[54] ));
 sky130_fd_sc_hd__dfrtp_1 _15305_ (.CLK(clknet_leaf_36_clk),
    .D(_00054_),
    .RESET_B(_00256_),
    .Q(\cycles[55] ));
 sky130_fd_sc_hd__dfrtp_1 _15306_ (.CLK(clknet_leaf_36_clk),
    .D(_00055_),
    .RESET_B(_00257_),
    .Q(\cycles[56] ));
 sky130_fd_sc_hd__dfrtp_1 _15307_ (.CLK(clknet_leaf_35_clk),
    .D(_00056_),
    .RESET_B(_00258_),
    .Q(\cycles[57] ));
 sky130_fd_sc_hd__dfrtp_1 _15308_ (.CLK(clknet_leaf_35_clk),
    .D(_00057_),
    .RESET_B(_00259_),
    .Q(\cycles[58] ));
 sky130_fd_sc_hd__dfrtp_1 _15309_ (.CLK(clknet_leaf_35_clk),
    .D(_00058_),
    .RESET_B(_00260_),
    .Q(\cycles[59] ));
 sky130_fd_sc_hd__dfrtp_1 _15310_ (.CLK(clknet_leaf_35_clk),
    .D(_00060_),
    .RESET_B(_00261_),
    .Q(\cycles[60] ));
 sky130_fd_sc_hd__dfrtp_1 _15311_ (.CLK(clknet_leaf_35_clk),
    .D(_00061_),
    .RESET_B(_00262_),
    .Q(\cycles[61] ));
 sky130_fd_sc_hd__dfrtp_1 _15312_ (.CLK(clknet_leaf_31_clk),
    .D(_00062_),
    .RESET_B(_00263_),
    .Q(\cycles[62] ));
 sky130_fd_sc_hd__dfrtp_1 _15313_ (.CLK(clknet_leaf_31_clk),
    .D(_00063_),
    .RESET_B(_00264_),
    .Q(\cycles[63] ));
 sky130_fd_sc_hd__dfrtp_2 _15314_ (.CLK(clknet_leaf_24_clk),
    .D(_01440_),
    .RESET_B(_00265_),
    .Q(\instr[0] ));
 sky130_fd_sc_hd__dfrtp_2 _15315_ (.CLK(clknet_leaf_24_clk),
    .D(_01441_),
    .RESET_B(_00266_),
    .Q(\instr[1] ));
 sky130_fd_sc_hd__dfrtp_2 _15316_ (.CLK(clknet_leaf_24_clk),
    .D(_01442_),
    .RESET_B(_00267_),
    .Q(\instr[2] ));
 sky130_fd_sc_hd__dfrtp_4 _15317_ (.CLK(clknet_leaf_24_clk),
    .D(_01443_),
    .RESET_B(_00268_),
    .Q(\instr[3] ));
 sky130_fd_sc_hd__dfrtp_1 _15318_ (.CLK(clknet_leaf_51_clk),
    .D(_01444_),
    .RESET_B(_00269_),
    .Q(\instr[4] ));
 sky130_fd_sc_hd__dfrtp_4 _15319_ (.CLK(clknet_leaf_24_clk),
    .D(_01445_),
    .RESET_B(_00270_),
    .Q(\instr[5] ));
 sky130_fd_sc_hd__dfrtp_2 _15320_ (.CLK(clknet_leaf_24_clk),
    .D(_01446_),
    .RESET_B(_00271_),
    .Q(\instr[6] ));
 sky130_fd_sc_hd__dfrtp_2 _15321_ (.CLK(clknet_leaf_52_clk),
    .D(_01447_),
    .RESET_B(_00272_),
    .Q(\B_type_imm[11] ));
 sky130_fd_sc_hd__dfrtp_4 _15322_ (.CLK(clknet_leaf_51_clk),
    .D(_01448_),
    .RESET_B(_00273_),
    .Q(\B_type_imm[1] ));
 sky130_fd_sc_hd__dfrtp_1 _15323_ (.CLK(clknet_leaf_50_clk),
    .D(_01449_),
    .RESET_B(_00274_),
    .Q(\B_type_imm[2] ));
 sky130_fd_sc_hd__dfrtp_1 _15324_ (.CLK(clknet_leaf_50_clk),
    .D(_01450_),
    .RESET_B(_00275_),
    .Q(\B_type_imm[3] ));
 sky130_fd_sc_hd__dfrtp_1 _15325_ (.CLK(clknet_leaf_50_clk),
    .D(_01451_),
    .RESET_B(_00276_),
    .Q(\B_type_imm[4] ));
 sky130_fd_sc_hd__dfrtp_4 _15326_ (.CLK(clknet_leaf_48_clk),
    .D(_01452_),
    .RESET_B(_00277_),
    .Q(\J_type_imm[12] ));
 sky130_fd_sc_hd__dfrtp_4 _15327_ (.CLK(clknet_leaf_52_clk),
    .D(_01453_),
    .RESET_B(_00278_),
    .Q(\J_type_imm[13] ));
 sky130_fd_sc_hd__dfrtp_4 _15328_ (.CLK(clknet_leaf_59_clk),
    .D(_01454_),
    .RESET_B(_00279_),
    .Q(\J_type_imm[14] ));
 sky130_fd_sc_hd__dfrtp_2 _15329_ (.CLK(clknet_leaf_57_clk),
    .D(_01455_),
    .RESET_B(_00280_),
    .Q(\J_type_imm[15] ));
 sky130_fd_sc_hd__dfrtp_1 _15330_ (.CLK(clknet_leaf_57_clk),
    .D(_01456_),
    .RESET_B(_00281_),
    .Q(\J_type_imm[16] ));
 sky130_fd_sc_hd__dfrtp_2 _15331_ (.CLK(clknet_leaf_53_clk),
    .D(_01457_),
    .RESET_B(_00282_),
    .Q(\J_type_imm[17] ));
 sky130_fd_sc_hd__dfrtp_2 _15332_ (.CLK(clknet_leaf_53_clk),
    .D(_01458_),
    .RESET_B(_00283_),
    .Q(\J_type_imm[18] ));
 sky130_fd_sc_hd__dfrtp_2 _15333_ (.CLK(clknet_leaf_57_clk),
    .D(_01459_),
    .RESET_B(_00284_),
    .Q(\J_type_imm[19] ));
 sky130_fd_sc_hd__dfrtp_2 _15334_ (.CLK(clknet_leaf_48_clk),
    .D(_01460_),
    .RESET_B(_00285_),
    .Q(\I_type_imm[0] ));
 sky130_fd_sc_hd__dfrtp_4 _15335_ (.CLK(clknet_leaf_52_clk),
    .D(_01461_),
    .RESET_B(_00286_),
    .Q(\I_type_imm[1] ));
 sky130_fd_sc_hd__dfrtp_2 _15336_ (.CLK(clknet_leaf_48_clk),
    .D(_01462_),
    .RESET_B(_00287_),
    .Q(\I_type_imm[2] ));
 sky130_fd_sc_hd__dfrtp_1 _15337_ (.CLK(clknet_leaf_48_clk),
    .D(_01463_),
    .RESET_B(_00288_),
    .Q(\I_type_imm[3] ));
 sky130_fd_sc_hd__dfrtp_1 _15338_ (.CLK(clknet_leaf_48_clk),
    .D(_01464_),
    .RESET_B(_00289_),
    .Q(\I_type_imm[4] ));
 sky130_fd_sc_hd__dfrtp_2 _15339_ (.CLK(clknet_leaf_42_clk),
    .D(_01465_),
    .RESET_B(_00290_),
    .Q(\B_type_imm[5] ));
 sky130_fd_sc_hd__dfrtp_2 _15340_ (.CLK(clknet_leaf_42_clk),
    .D(_01466_),
    .RESET_B(_00291_),
    .Q(\B_type_imm[6] ));
 sky130_fd_sc_hd__dfrtp_2 _15341_ (.CLK(clknet_leaf_43_clk),
    .D(_01467_),
    .RESET_B(_00292_),
    .Q(\B_type_imm[7] ));
 sky130_fd_sc_hd__dfrtp_2 _15342_ (.CLK(clknet_leaf_49_clk),
    .D(_01468_),
    .RESET_B(_00293_),
    .Q(\B_type_imm[8] ));
 sky130_fd_sc_hd__dfrtp_1 _15343_ (.CLK(clknet_leaf_49_clk),
    .D(_01469_),
    .RESET_B(_00294_),
    .Q(\B_type_imm[9] ));
 sky130_fd_sc_hd__dfrtp_4 _15344_ (.CLK(clknet_leaf_49_clk),
    .D(_01470_),
    .RESET_B(_00295_),
    .Q(\barrel_shifter_right.arith ));
 sky130_fd_sc_hd__dfrtp_4 _15345_ (.CLK(clknet_leaf_47_clk),
    .D(_01471_),
    .RESET_B(_00296_),
    .Q(\B_type_imm[12] ));
 sky130_fd_sc_hd__dfxtp_1 _15346_ (.CLK(clknet_leaf_120_clk),
    .D(_01472_),
    .Q(\regs[17][0] ));
 sky130_fd_sc_hd__dfxtp_1 _15347_ (.CLK(clknet_leaf_132_clk),
    .D(_01473_),
    .Q(\regs[17][1] ));
 sky130_fd_sc_hd__dfxtp_1 _15348_ (.CLK(clknet_leaf_132_clk),
    .D(_01474_),
    .Q(\regs[17][2] ));
 sky130_fd_sc_hd__dfxtp_1 _15349_ (.CLK(clknet_leaf_4_clk),
    .D(_01475_),
    .Q(\regs[17][3] ));
 sky130_fd_sc_hd__dfxtp_1 _15350_ (.CLK(clknet_leaf_122_clk),
    .D(_01476_),
    .Q(\regs[17][4] ));
 sky130_fd_sc_hd__dfxtp_1 _15351_ (.CLK(clknet_leaf_4_clk),
    .D(_01477_),
    .Q(\regs[17][5] ));
 sky130_fd_sc_hd__dfxtp_1 _15352_ (.CLK(clknet_leaf_108_clk),
    .D(_01478_),
    .Q(\regs[17][6] ));
 sky130_fd_sc_hd__dfxtp_1 _15353_ (.CLK(clknet_leaf_123_clk),
    .D(_01479_),
    .Q(\regs[17][7] ));
 sky130_fd_sc_hd__dfxtp_1 _15354_ (.CLK(clknet_leaf_4_clk),
    .D(_01480_),
    .Q(\regs[17][8] ));
 sky130_fd_sc_hd__dfxtp_1 _15355_ (.CLK(clknet_leaf_124_clk),
    .D(_01481_),
    .Q(\regs[17][9] ));
 sky130_fd_sc_hd__dfxtp_1 _15356_ (.CLK(clknet_leaf_70_clk),
    .D(_01482_),
    .Q(\regs[17][10] ));
 sky130_fd_sc_hd__dfxtp_1 _15357_ (.CLK(clknet_leaf_86_clk),
    .D(_01483_),
    .Q(\regs[17][11] ));
 sky130_fd_sc_hd__dfxtp_1 _15358_ (.CLK(clknet_leaf_87_clk),
    .D(_01484_),
    .Q(\regs[17][12] ));
 sky130_fd_sc_hd__dfxtp_1 _15359_ (.CLK(clknet_leaf_86_clk),
    .D(_01485_),
    .Q(\regs[17][13] ));
 sky130_fd_sc_hd__dfxtp_1 _15360_ (.CLK(clknet_leaf_83_clk),
    .D(_01486_),
    .Q(\regs[17][14] ));
 sky130_fd_sc_hd__dfxtp_1 _15361_ (.CLK(clknet_leaf_112_clk),
    .D(_01487_),
    .Q(\regs[17][15] ));
 sky130_fd_sc_hd__dfxtp_1 _15362_ (.CLK(clknet_leaf_82_clk),
    .D(_01488_),
    .Q(\regs[17][16] ));
 sky130_fd_sc_hd__dfxtp_1 _15363_ (.CLK(clknet_leaf_65_clk),
    .D(_01489_),
    .Q(\regs[17][17] ));
 sky130_fd_sc_hd__dfxtp_1 _15364_ (.CLK(clknet_leaf_74_clk),
    .D(_01490_),
    .Q(\regs[17][18] ));
 sky130_fd_sc_hd__dfxtp_1 _15365_ (.CLK(clknet_leaf_84_clk),
    .D(_01491_),
    .Q(\regs[17][19] ));
 sky130_fd_sc_hd__dfxtp_1 _15366_ (.CLK(clknet_leaf_26_clk),
    .D(_01492_),
    .Q(\regs[17][20] ));
 sky130_fd_sc_hd__dfxtp_1 _15367_ (.CLK(clknet_leaf_51_clk),
    .D(_01493_),
    .Q(\regs[17][21] ));
 sky130_fd_sc_hd__dfxtp_1 _15368_ (.CLK(clknet_leaf_53_clk),
    .D(_01494_),
    .Q(\regs[17][22] ));
 sky130_fd_sc_hd__dfxtp_1 _15369_ (.CLK(clknet_leaf_25_clk),
    .D(_01495_),
    .Q(\regs[17][23] ));
 sky130_fd_sc_hd__dfxtp_1 _15370_ (.CLK(clknet_leaf_23_clk),
    .D(_01496_),
    .Q(\regs[17][24] ));
 sky130_fd_sc_hd__dfxtp_1 _15371_ (.CLK(clknet_leaf_21_clk),
    .D(_01497_),
    .Q(\regs[17][25] ));
 sky130_fd_sc_hd__dfxtp_1 _15372_ (.CLK(clknet_leaf_53_clk),
    .D(_01498_),
    .Q(\regs[17][26] ));
 sky130_fd_sc_hd__dfxtp_1 _15373_ (.CLK(clknet_leaf_57_clk),
    .D(_01499_),
    .Q(\regs[17][27] ));
 sky130_fd_sc_hd__dfxtp_1 _15374_ (.CLK(clknet_leaf_26_clk),
    .D(_01500_),
    .Q(\regs[17][28] ));
 sky130_fd_sc_hd__dfxtp_1 _15375_ (.CLK(clknet_leaf_51_clk),
    .D(_01501_),
    .Q(\regs[17][29] ));
 sky130_fd_sc_hd__dfxtp_1 _15376_ (.CLK(clknet_leaf_55_clk),
    .D(_01502_),
    .Q(\regs[17][30] ));
 sky130_fd_sc_hd__dfxtp_1 _15377_ (.CLK(clknet_leaf_71_clk),
    .D(_01503_),
    .Q(\regs[17][31] ));
 sky130_fd_sc_hd__dfrtp_1 _15378_ (.CLK(clknet_leaf_50_clk),
    .D(_01504_),
    .RESET_B(_00297_),
    .Q(\PC[2] ));
 sky130_fd_sc_hd__dfrtp_4 _15379_ (.CLK(clknet_leaf_42_clk),
    .D(_01505_),
    .RESET_B(_00298_),
    .Q(\PC[3] ));
 sky130_fd_sc_hd__dfrtp_4 _15380_ (.CLK(clknet_leaf_43_clk),
    .D(_01506_),
    .RESET_B(_00299_),
    .Q(\PC[4] ));
 sky130_fd_sc_hd__dfrtp_2 _15381_ (.CLK(clknet_leaf_43_clk),
    .D(_01507_),
    .RESET_B(_00300_),
    .Q(\PC[5] ));
 sky130_fd_sc_hd__dfrtp_1 _15382_ (.CLK(clknet_leaf_44_clk),
    .D(_01508_),
    .RESET_B(_00301_),
    .Q(\PC[6] ));
 sky130_fd_sc_hd__dfrtp_4 _15383_ (.CLK(clknet_leaf_44_clk),
    .D(_01509_),
    .RESET_B(_00302_),
    .Q(\PC[7] ));
 sky130_fd_sc_hd__dfrtp_2 _15384_ (.CLK(clknet_leaf_45_clk),
    .D(_01510_),
    .RESET_B(_00303_),
    .Q(\PC[8] ));
 sky130_fd_sc_hd__dfrtp_4 _15385_ (.CLK(clknet_leaf_45_clk),
    .D(_01511_),
    .RESET_B(_00304_),
    .Q(\PC[9] ));
 sky130_fd_sc_hd__dfrtp_2 _15386_ (.CLK(clknet_leaf_45_clk),
    .D(_01512_),
    .RESET_B(_00305_),
    .Q(\PC[10] ));
 sky130_fd_sc_hd__dfrtp_4 _15387_ (.CLK(clknet_leaf_45_clk),
    .D(_01513_),
    .RESET_B(_00306_),
    .Q(\PC[11] ));
 sky130_fd_sc_hd__dfrtp_1 _15388_ (.CLK(clknet_leaf_47_clk),
    .D(_01514_),
    .RESET_B(_00307_),
    .Q(\PC[12] ));
 sky130_fd_sc_hd__dfrtp_4 _15389_ (.CLK(clknet_leaf_46_clk),
    .D(_01515_),
    .RESET_B(_00308_),
    .Q(\PC[13] ));
 sky130_fd_sc_hd__dfrtp_4 _15390_ (.CLK(clknet_leaf_60_clk),
    .D(_01516_),
    .RESET_B(_00309_),
    .Q(\PC[14] ));
 sky130_fd_sc_hd__dfrtp_1 _15391_ (.CLK(clknet_leaf_59_clk),
    .D(_01517_),
    .RESET_B(_00310_),
    .Q(\PC[15] ));
 sky130_fd_sc_hd__dfrtp_4 _15392_ (.CLK(clknet_leaf_60_clk),
    .D(_01518_),
    .RESET_B(_00311_),
    .Q(\PC[16] ));
 sky130_fd_sc_hd__dfrtp_4 _15393_ (.CLK(clknet_leaf_61_clk),
    .D(_01519_),
    .RESET_B(_00312_),
    .Q(\PC[17] ));
 sky130_fd_sc_hd__dfrtp_4 _15394_ (.CLK(clknet_leaf_60_clk),
    .D(_01520_),
    .RESET_B(_00313_),
    .Q(\PC[18] ));
 sky130_fd_sc_hd__dfrtp_4 _15395_ (.CLK(clknet_leaf_46_clk),
    .D(_01521_),
    .RESET_B(_00314_),
    .Q(\PC[19] ));
 sky130_fd_sc_hd__dfrtp_1 _15396_ (.CLK(clknet_leaf_45_clk),
    .D(_01522_),
    .RESET_B(_00315_),
    .Q(\PC[20] ));
 sky130_fd_sc_hd__dfrtp_4 _15397_ (.CLK(clknet_leaf_45_clk),
    .D(_01523_),
    .RESET_B(_00316_),
    .Q(\PC[21] ));
 sky130_fd_sc_hd__dfrtp_4 _15398_ (.CLK(clknet_leaf_61_clk),
    .D(_01524_),
    .RESET_B(_00317_),
    .Q(\PC[22] ));
 sky130_fd_sc_hd__dfrtp_4 _15399_ (.CLK(clknet_leaf_61_clk),
    .D(_01525_),
    .RESET_B(_00318_),
    .Q(\PC[23] ));
 sky130_fd_sc_hd__conb_1 leorv32_99 (.LO(net99));
 sky130_fd_sc_hd__conb_1 leorv32_100 (.LO(net100));
 sky130_fd_sc_hd__conb_1 leorv32_101 (.LO(net101));
 sky130_fd_sc_hd__conb_1 leorv32_102 (.LO(net102));
 sky130_fd_sc_hd__conb_1 leorv32_103 (.LO(net103));
 sky130_fd_sc_hd__conb_1 leorv32_104 (.LO(net104));
 sky130_fd_sc_hd__conb_1 leorv32_105 (.LO(net105));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_0_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_0_clk));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__decap_3 PHY_204 ();
 sky130_fd_sc_hd__decap_3 PHY_205 ();
 sky130_fd_sc_hd__decap_3 PHY_206 ();
 sky130_fd_sc_hd__decap_3 PHY_207 ();
 sky130_fd_sc_hd__decap_3 PHY_208 ();
 sky130_fd_sc_hd__decap_3 PHY_209 ();
 sky130_fd_sc_hd__decap_3 PHY_210 ();
 sky130_fd_sc_hd__decap_3 PHY_211 ();
 sky130_fd_sc_hd__decap_3 PHY_212 ();
 sky130_fd_sc_hd__decap_3 PHY_213 ();
 sky130_fd_sc_hd__decap_3 PHY_214 ();
 sky130_fd_sc_hd__decap_3 PHY_215 ();
 sky130_fd_sc_hd__decap_3 PHY_216 ();
 sky130_fd_sc_hd__decap_3 PHY_217 ();
 sky130_fd_sc_hd__decap_3 PHY_218 ();
 sky130_fd_sc_hd__decap_3 PHY_219 ();
 sky130_fd_sc_hd__decap_3 PHY_220 ();
 sky130_fd_sc_hd__decap_3 PHY_221 ();
 sky130_fd_sc_hd__decap_3 PHY_222 ();
 sky130_fd_sc_hd__decap_3 PHY_223 ();
 sky130_fd_sc_hd__decap_3 PHY_224 ();
 sky130_fd_sc_hd__decap_3 PHY_225 ();
 sky130_fd_sc_hd__decap_3 PHY_226 ();
 sky130_fd_sc_hd__decap_3 PHY_227 ();
 sky130_fd_sc_hd__decap_3 PHY_228 ();
 sky130_fd_sc_hd__decap_3 PHY_229 ();
 sky130_fd_sc_hd__decap_3 PHY_230 ();
 sky130_fd_sc_hd__decap_3 PHY_231 ();
 sky130_fd_sc_hd__decap_3 PHY_232 ();
 sky130_fd_sc_hd__decap_3 PHY_233 ();
 sky130_fd_sc_hd__decap_3 PHY_234 ();
 sky130_fd_sc_hd__decap_3 PHY_235 ();
 sky130_fd_sc_hd__decap_3 PHY_236 ();
 sky130_fd_sc_hd__decap_3 PHY_237 ();
 sky130_fd_sc_hd__decap_3 PHY_238 ();
 sky130_fd_sc_hd__decap_3 PHY_239 ();
 sky130_fd_sc_hd__decap_3 PHY_240 ();
 sky130_fd_sc_hd__decap_3 PHY_241 ();
 sky130_fd_sc_hd__decap_3 PHY_242 ();
 sky130_fd_sc_hd__decap_3 PHY_243 ();
 sky130_fd_sc_hd__decap_3 PHY_244 ();
 sky130_fd_sc_hd__decap_3 PHY_245 ();
 sky130_fd_sc_hd__decap_3 PHY_246 ();
 sky130_fd_sc_hd__decap_3 PHY_247 ();
 sky130_fd_sc_hd__decap_3 PHY_248 ();
 sky130_fd_sc_hd__decap_3 PHY_249 ();
 sky130_fd_sc_hd__decap_3 PHY_250 ();
 sky130_fd_sc_hd__decap_3 PHY_251 ();
 sky130_fd_sc_hd__decap_3 PHY_252 ();
 sky130_fd_sc_hd__decap_3 PHY_253 ();
 sky130_fd_sc_hd__decap_3 PHY_254 ();
 sky130_fd_sc_hd__decap_3 PHY_255 ();
 sky130_fd_sc_hd__decap_3 PHY_256 ();
 sky130_fd_sc_hd__decap_3 PHY_257 ();
 sky130_fd_sc_hd__decap_3 PHY_258 ();
 sky130_fd_sc_hd__decap_3 PHY_259 ();
 sky130_fd_sc_hd__decap_3 PHY_260 ();
 sky130_fd_sc_hd__decap_3 PHY_261 ();
 sky130_fd_sc_hd__decap_3 PHY_262 ();
 sky130_fd_sc_hd__decap_3 PHY_263 ();
 sky130_fd_sc_hd__decap_3 PHY_264 ();
 sky130_fd_sc_hd__decap_3 PHY_265 ();
 sky130_fd_sc_hd__decap_3 PHY_266 ();
 sky130_fd_sc_hd__decap_3 PHY_267 ();
 sky130_fd_sc_hd__decap_3 PHY_268 ();
 sky130_fd_sc_hd__decap_3 PHY_269 ();
 sky130_fd_sc_hd__decap_3 PHY_270 ();
 sky130_fd_sc_hd__decap_3 PHY_271 ();
 sky130_fd_sc_hd__decap_3 PHY_272 ();
 sky130_fd_sc_hd__decap_3 PHY_273 ();
 sky130_fd_sc_hd__decap_3 PHY_274 ();
 sky130_fd_sc_hd__decap_3 PHY_275 ();
 sky130_fd_sc_hd__decap_3 PHY_276 ();
 sky130_fd_sc_hd__decap_3 PHY_277 ();
 sky130_fd_sc_hd__decap_3 PHY_278 ();
 sky130_fd_sc_hd__decap_3 PHY_279 ();
 sky130_fd_sc_hd__decap_3 PHY_280 ();
 sky130_fd_sc_hd__decap_3 PHY_281 ();
 sky130_fd_sc_hd__decap_3 PHY_282 ();
 sky130_fd_sc_hd__decap_3 PHY_283 ();
 sky130_fd_sc_hd__decap_3 PHY_284 ();
 sky130_fd_sc_hd__decap_3 PHY_285 ();
 sky130_fd_sc_hd__decap_3 PHY_286 ();
 sky130_fd_sc_hd__decap_3 PHY_287 ();
 sky130_fd_sc_hd__decap_3 PHY_288 ();
 sky130_fd_sc_hd__decap_3 PHY_289 ();
 sky130_fd_sc_hd__decap_3 PHY_290 ();
 sky130_fd_sc_hd__decap_3 PHY_291 ();
 sky130_fd_sc_hd__decap_3 PHY_292 ();
 sky130_fd_sc_hd__decap_3 PHY_293 ();
 sky130_fd_sc_hd__decap_3 PHY_294 ();
 sky130_fd_sc_hd__decap_3 PHY_295 ();
 sky130_fd_sc_hd__decap_3 PHY_296 ();
 sky130_fd_sc_hd__decap_3 PHY_297 ();
 sky130_fd_sc_hd__decap_3 PHY_298 ();
 sky130_fd_sc_hd__decap_3 PHY_299 ();
 sky130_fd_sc_hd__decap_3 PHY_300 ();
 sky130_fd_sc_hd__decap_3 PHY_301 ();
 sky130_fd_sc_hd__decap_3 PHY_302 ();
 sky130_fd_sc_hd__decap_3 PHY_303 ();
 sky130_fd_sc_hd__decap_3 PHY_304 ();
 sky130_fd_sc_hd__decap_3 PHY_305 ();
 sky130_fd_sc_hd__decap_3 PHY_306 ();
 sky130_fd_sc_hd__decap_3 PHY_307 ();
 sky130_fd_sc_hd__decap_3 PHY_308 ();
 sky130_fd_sc_hd__decap_3 PHY_309 ();
 sky130_fd_sc_hd__decap_3 PHY_310 ();
 sky130_fd_sc_hd__decap_3 PHY_311 ();
 sky130_fd_sc_hd__decap_3 PHY_312 ();
 sky130_fd_sc_hd__decap_3 PHY_313 ();
 sky130_fd_sc_hd__decap_3 PHY_314 ();
 sky130_fd_sc_hd__decap_3 PHY_315 ();
 sky130_fd_sc_hd__decap_3 PHY_316 ();
 sky130_fd_sc_hd__decap_3 PHY_317 ();
 sky130_fd_sc_hd__decap_3 PHY_318 ();
 sky130_fd_sc_hd__decap_3 PHY_319 ();
 sky130_fd_sc_hd__decap_3 PHY_320 ();
 sky130_fd_sc_hd__decap_3 PHY_321 ();
 sky130_fd_sc_hd__decap_3 PHY_322 ();
 sky130_fd_sc_hd__decap_3 PHY_323 ();
 sky130_fd_sc_hd__decap_3 PHY_324 ();
 sky130_fd_sc_hd__decap_3 PHY_325 ();
 sky130_fd_sc_hd__decap_3 PHY_326 ();
 sky130_fd_sc_hd__decap_3 PHY_327 ();
 sky130_fd_sc_hd__decap_3 PHY_328 ();
 sky130_fd_sc_hd__decap_3 PHY_329 ();
 sky130_fd_sc_hd__decap_3 PHY_330 ();
 sky130_fd_sc_hd__decap_3 PHY_331 ();
 sky130_fd_sc_hd__decap_3 PHY_332 ();
 sky130_fd_sc_hd__decap_3 PHY_333 ();
 sky130_fd_sc_hd__decap_3 PHY_334 ();
 sky130_fd_sc_hd__decap_3 PHY_335 ();
 sky130_fd_sc_hd__decap_3 PHY_336 ();
 sky130_fd_sc_hd__decap_3 PHY_337 ();
 sky130_fd_sc_hd__decap_3 PHY_338 ();
 sky130_fd_sc_hd__decap_3 PHY_339 ();
 sky130_fd_sc_hd__decap_3 PHY_340 ();
 sky130_fd_sc_hd__decap_3 PHY_341 ();
 sky130_fd_sc_hd__decap_3 PHY_342 ();
 sky130_fd_sc_hd__decap_3 PHY_343 ();
 sky130_fd_sc_hd__decap_3 PHY_344 ();
 sky130_fd_sc_hd__decap_3 PHY_345 ();
 sky130_fd_sc_hd__decap_3 PHY_346 ();
 sky130_fd_sc_hd__decap_3 PHY_347 ();
 sky130_fd_sc_hd__decap_3 PHY_348 ();
 sky130_fd_sc_hd__decap_3 PHY_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3623 ();
 sky130_fd_sc_hd__buf_4 input1 (.A(mem_rbusy),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_4 input2 (.A(mem_rdata[0]),
    .X(net2));
 sky130_fd_sc_hd__buf_2 input3 (.A(mem_rdata[10]),
    .X(net3));
 sky130_fd_sc_hd__buf_2 input4 (.A(mem_rdata[11]),
    .X(net4));
 sky130_fd_sc_hd__buf_2 input5 (.A(mem_rdata[12]),
    .X(net5));
 sky130_fd_sc_hd__buf_2 input6 (.A(mem_rdata[13]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_4 input7 (.A(mem_rdata[14]),
    .X(net7));
 sky130_fd_sc_hd__buf_4 input8 (.A(mem_rdata[15]),
    .X(net8));
 sky130_fd_sc_hd__buf_4 input9 (.A(mem_rdata[16]),
    .X(net9));
 sky130_fd_sc_hd__buf_6 input10 (.A(mem_rdata[17]),
    .X(net10));
 sky130_fd_sc_hd__buf_4 input11 (.A(mem_rdata[18]),
    .X(net11));
 sky130_fd_sc_hd__buf_8 input12 (.A(mem_rdata[19]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_4 input13 (.A(mem_rdata[1]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_4 input14 (.A(mem_rdata[20]),
    .X(net14));
 sky130_fd_sc_hd__buf_6 input15 (.A(mem_rdata[21]),
    .X(net15));
 sky130_fd_sc_hd__buf_8 input16 (.A(mem_rdata[22]),
    .X(net16));
 sky130_fd_sc_hd__buf_4 input17 (.A(mem_rdata[23]),
    .X(net17));
 sky130_fd_sc_hd__buf_8 input18 (.A(mem_rdata[24]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_2 input19 (.A(mem_rdata[25]),
    .X(net19));
 sky130_fd_sc_hd__buf_2 input20 (.A(mem_rdata[26]),
    .X(net20));
 sky130_fd_sc_hd__buf_2 input21 (.A(mem_rdata[27]),
    .X(net21));
 sky130_fd_sc_hd__buf_2 input22 (.A(mem_rdata[28]),
    .X(net22));
 sky130_fd_sc_hd__buf_2 input23 (.A(mem_rdata[29]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_4 input24 (.A(mem_rdata[2]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_4 input25 (.A(mem_rdata[30]),
    .X(net25));
 sky130_fd_sc_hd__buf_2 input26 (.A(mem_rdata[31]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_4 input27 (.A(mem_rdata[3]),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_4 input28 (.A(mem_rdata[4]),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_4 input29 (.A(mem_rdata[5]),
    .X(net29));
 sky130_fd_sc_hd__buf_2 input30 (.A(mem_rdata[6]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_4 input31 (.A(mem_rdata[7]),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_4 input32 (.A(mem_rdata[8]),
    .X(net32));
 sky130_fd_sc_hd__buf_2 input33 (.A(mem_rdata[9]),
    .X(net33));
 sky130_fd_sc_hd__buf_4 input34 (.A(mem_wbusy),
    .X(net34));
 sky130_fd_sc_hd__buf_2 input35 (.A(mhartid_0),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_1 input36 (.A(reset),
    .X(net36));
 sky130_fd_sc_hd__buf_2 output37 (.A(net37),
    .X(mem_addr[0]));
 sky130_fd_sc_hd__buf_2 output38 (.A(net38),
    .X(mem_addr[10]));
 sky130_fd_sc_hd__buf_2 output39 (.A(net39),
    .X(mem_addr[11]));
 sky130_fd_sc_hd__buf_2 output40 (.A(net40),
    .X(mem_addr[12]));
 sky130_fd_sc_hd__buf_2 output41 (.A(net41),
    .X(mem_addr[13]));
 sky130_fd_sc_hd__buf_2 output42 (.A(net42),
    .X(mem_addr[14]));
 sky130_fd_sc_hd__buf_2 output43 (.A(net43),
    .X(mem_addr[15]));
 sky130_fd_sc_hd__buf_2 output44 (.A(net44),
    .X(mem_addr[16]));
 sky130_fd_sc_hd__buf_2 output45 (.A(net45),
    .X(mem_addr[17]));
 sky130_fd_sc_hd__buf_2 output46 (.A(net46),
    .X(mem_addr[18]));
 sky130_fd_sc_hd__buf_2 output47 (.A(net47),
    .X(mem_addr[19]));
 sky130_fd_sc_hd__buf_2 output48 (.A(net48),
    .X(mem_addr[1]));
 sky130_fd_sc_hd__buf_2 output49 (.A(net49),
    .X(mem_addr[20]));
 sky130_fd_sc_hd__buf_2 output50 (.A(net50),
    .X(mem_addr[21]));
 sky130_fd_sc_hd__buf_2 output51 (.A(net51),
    .X(mem_addr[22]));
 sky130_fd_sc_hd__buf_2 output52 (.A(net52),
    .X(mem_addr[23]));
 sky130_fd_sc_hd__buf_2 output53 (.A(net53),
    .X(mem_addr[2]));
 sky130_fd_sc_hd__buf_2 output54 (.A(net54),
    .X(mem_addr[3]));
 sky130_fd_sc_hd__buf_2 output55 (.A(net55),
    .X(mem_addr[4]));
 sky130_fd_sc_hd__buf_2 output56 (.A(net56),
    .X(mem_addr[5]));
 sky130_fd_sc_hd__buf_2 output57 (.A(net57),
    .X(mem_addr[6]));
 sky130_fd_sc_hd__buf_2 output58 (.A(net58),
    .X(mem_addr[7]));
 sky130_fd_sc_hd__buf_2 output59 (.A(net59),
    .X(mem_addr[8]));
 sky130_fd_sc_hd__buf_2 output60 (.A(net60),
    .X(mem_addr[9]));
 sky130_fd_sc_hd__buf_2 output61 (.A(net61),
    .X(mem_rstrb));
 sky130_fd_sc_hd__buf_2 output62 (.A(net62),
    .X(mem_wdata[0]));
 sky130_fd_sc_hd__buf_2 output63 (.A(net63),
    .X(mem_wdata[10]));
 sky130_fd_sc_hd__buf_2 output64 (.A(net64),
    .X(mem_wdata[11]));
 sky130_fd_sc_hd__buf_2 output65 (.A(net65),
    .X(mem_wdata[12]));
 sky130_fd_sc_hd__buf_2 output66 (.A(net66),
    .X(mem_wdata[13]));
 sky130_fd_sc_hd__buf_2 output67 (.A(net67),
    .X(mem_wdata[14]));
 sky130_fd_sc_hd__buf_2 output68 (.A(net68),
    .X(mem_wdata[15]));
 sky130_fd_sc_hd__buf_2 output69 (.A(net69),
    .X(mem_wdata[16]));
 sky130_fd_sc_hd__buf_2 output70 (.A(net70),
    .X(mem_wdata[17]));
 sky130_fd_sc_hd__buf_2 output71 (.A(net71),
    .X(mem_wdata[18]));
 sky130_fd_sc_hd__buf_2 output72 (.A(net72),
    .X(mem_wdata[19]));
 sky130_fd_sc_hd__buf_2 output73 (.A(net73),
    .X(mem_wdata[1]));
 sky130_fd_sc_hd__buf_2 output74 (.A(net74),
    .X(mem_wdata[20]));
 sky130_fd_sc_hd__buf_2 output75 (.A(net75),
    .X(mem_wdata[21]));
 sky130_fd_sc_hd__buf_2 output76 (.A(net76),
    .X(mem_wdata[22]));
 sky130_fd_sc_hd__buf_2 output77 (.A(net77),
    .X(mem_wdata[23]));
 sky130_fd_sc_hd__buf_2 output78 (.A(net78),
    .X(mem_wdata[24]));
 sky130_fd_sc_hd__buf_2 output79 (.A(net79),
    .X(mem_wdata[25]));
 sky130_fd_sc_hd__buf_2 output80 (.A(net80),
    .X(mem_wdata[26]));
 sky130_fd_sc_hd__buf_2 output81 (.A(net81),
    .X(mem_wdata[27]));
 sky130_fd_sc_hd__buf_2 output82 (.A(net82),
    .X(mem_wdata[28]));
 sky130_fd_sc_hd__buf_2 output83 (.A(net83),
    .X(mem_wdata[29]));
 sky130_fd_sc_hd__buf_2 output84 (.A(net84),
    .X(mem_wdata[2]));
 sky130_fd_sc_hd__buf_2 output85 (.A(net85),
    .X(mem_wdata[30]));
 sky130_fd_sc_hd__buf_2 output86 (.A(net86),
    .X(mem_wdata[31]));
 sky130_fd_sc_hd__buf_2 output87 (.A(net87),
    .X(mem_wdata[3]));
 sky130_fd_sc_hd__buf_2 output88 (.A(net88),
    .X(mem_wdata[4]));
 sky130_fd_sc_hd__buf_2 output89 (.A(net89),
    .X(mem_wdata[5]));
 sky130_fd_sc_hd__buf_2 output90 (.A(net90),
    .X(mem_wdata[6]));
 sky130_fd_sc_hd__buf_2 output91 (.A(net91),
    .X(mem_wdata[7]));
 sky130_fd_sc_hd__buf_2 output92 (.A(net92),
    .X(mem_wdata[8]));
 sky130_fd_sc_hd__buf_2 output93 (.A(net93),
    .X(mem_wdata[9]));
 sky130_fd_sc_hd__buf_2 output94 (.A(net94),
    .X(mem_wmask[0]));
 sky130_fd_sc_hd__buf_2 output95 (.A(net95),
    .X(mem_wmask[1]));
 sky130_fd_sc_hd__buf_2 output96 (.A(net96),
    .X(mem_wmask[2]));
 sky130_fd_sc_hd__buf_2 output97 (.A(net97),
    .X(mem_wmask[3]));
 sky130_fd_sc_hd__conb_1 leorv32_98 (.LO(net98));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_1_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_1_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_2_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_2_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_3_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_3_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_4_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_4_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_5_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_5_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_6_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_6_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_7_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_7_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_8_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_8_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_9_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_9_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_10_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_10_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_11_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_11_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_12_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_12_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_13_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_13_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_14_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_14_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_15_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_15_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_16_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_16_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_17_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_17_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_18_clk (.A(clknet_opt_3_0_clk),
    .X(clknet_leaf_18_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_19_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_19_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_20_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_20_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_21_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_21_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_22_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_22_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_23_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_23_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_24_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_24_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_25_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_25_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_26_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_26_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_27_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_27_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_28_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_28_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_29_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_29_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_30_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_30_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_31_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_31_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_32_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_32_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_33_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_33_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_34_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_34_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_35_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_35_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_36_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_36_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_37_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_37_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_38_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_38_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_39_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_39_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_40_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_40_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_41_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_41_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_42_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_42_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_43_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_43_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_44_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_44_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_45_clk (.A(clknet_opt_2_0_clk),
    .X(clknet_leaf_45_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_46_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_46_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_47_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_47_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_48_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_48_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_49_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_49_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_50_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_50_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_51_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_51_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_52_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_52_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_53_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_53_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_54_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_54_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_55_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_55_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_56_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_56_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_57_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_57_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_59_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_59_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_60_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_60_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_61_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_61_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_62_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_62_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_63_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_63_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_64_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_64_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_65_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_65_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_66_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_66_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_67_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_67_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_68_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_68_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_69_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_69_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_70_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_70_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_71_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_71_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_72_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_72_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_73_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_73_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_74_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_74_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_75_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_75_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_76_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_76_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_77_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_77_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_78_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_78_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_79_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_79_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_80_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_80_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_81_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_81_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_82_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_82_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_83_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_83_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_84_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_84_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_85_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_85_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_86_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_86_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_87_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_87_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_88_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_88_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_89_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_89_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_90_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_90_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_91_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_91_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_92_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_92_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_93_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_93_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_94_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_94_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_95_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_95_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_96_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_96_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_97_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_97_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_98_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_98_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_99_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_99_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_100_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_100_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_101_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_101_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_102_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_102_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_103_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_103_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_104_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_104_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_105_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_105_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_106_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_106_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_107_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_107_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_108_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_108_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_109_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_109_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_110_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_110_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_111_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_111_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_112_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_112_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_113_clk (.A(clknet_opt_1_0_clk),
    .X(clknet_leaf_113_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_114_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_114_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_115_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_115_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_116_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_116_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_117_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_117_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_118_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_118_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_119_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_119_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_120_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_120_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_121_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_121_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_122_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_122_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_123_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_123_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_124_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_124_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_125_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_125_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_126_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_126_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_127_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_127_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_128_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_128_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_129_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_129_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_130_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_130_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_131_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_131_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_132_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_132_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_133_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_133_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_134_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_134_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_135_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_135_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_1_0_0_clk (.A(clknet_0_clk),
    .X(clknet_1_0_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_1_1_0_clk (.A(clknet_0_clk),
    .X(clknet_1_1_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_0_0_clk (.A(clknet_1_0_0_clk),
    .X(clknet_2_0_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_1_0_clk (.A(clknet_1_0_0_clk),
    .X(clknet_2_1_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_2_0_clk (.A(clknet_1_1_0_clk),
    .X(clknet_2_2_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_3_0_clk (.A(clknet_1_1_0_clk),
    .X(clknet_2_3_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_0_0_clk (.A(clknet_2_0_0_clk),
    .X(clknet_3_0_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_1_0_clk (.A(clknet_2_0_0_clk),
    .X(clknet_3_1_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_2_0_clk (.A(clknet_2_1_0_clk),
    .X(clknet_3_2_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_3_0_clk (.A(clknet_2_1_0_clk),
    .X(clknet_3_3_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_4_0_clk (.A(clknet_2_2_0_clk),
    .X(clknet_3_4_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_5_0_clk (.A(clknet_2_2_0_clk),
    .X(clknet_3_5_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_6_0_clk (.A(clknet_2_3_0_clk),
    .X(clknet_3_6_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_7_0_clk (.A(clknet_2_3_0_clk),
    .X(clknet_3_7_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_0_0_clk (.A(clknet_3_0_0_clk),
    .X(clknet_4_0_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_1_0_clk (.A(clknet_3_0_0_clk),
    .X(clknet_4_1_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_2_0_clk (.A(clknet_3_1_0_clk),
    .X(clknet_4_2_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_3_0_clk (.A(clknet_3_1_0_clk),
    .X(clknet_4_3_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_4_0_clk (.A(clknet_3_2_0_clk),
    .X(clknet_4_4_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_5_0_clk (.A(clknet_3_2_0_clk),
    .X(clknet_4_5_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_6_0_clk (.A(clknet_3_3_0_clk),
    .X(clknet_4_6_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_7_0_clk (.A(clknet_3_3_0_clk),
    .X(clknet_4_7_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_8_0_clk (.A(clknet_3_4_0_clk),
    .X(clknet_4_8_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_9_0_clk (.A(clknet_3_4_0_clk),
    .X(clknet_4_9_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_10_0_clk (.A(clknet_3_5_0_clk),
    .X(clknet_4_10_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_11_0_clk (.A(clknet_3_5_0_clk),
    .X(clknet_4_11_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_12_0_clk (.A(clknet_3_6_0_clk),
    .X(clknet_4_12_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_13_0_clk (.A(clknet_3_6_0_clk),
    .X(clknet_4_13_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_14_0_clk (.A(clknet_3_7_0_clk),
    .X(clknet_4_14_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_15_0_clk (.A(clknet_3_7_0_clk),
    .X(clknet_4_15_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_1_0_clk (.A(clknet_4_4_0_clk),
    .X(clknet_opt_1_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_2_0_clk (.A(clknet_4_11_0_clk),
    .X(clknet_opt_2_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_3_0_clk (.A(clknet_4_12_0_clk),
    .X(clknet_opt_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__10269__B1 (.DIODE(\B_type_imm[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10195__A (.DIODE(\B_type_imm[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07441__A (.DIODE(\B_type_imm[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07438__A (.DIODE(\B_type_imm[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07435__A (.DIODE(\B_type_imm[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07434__A (.DIODE(\B_type_imm[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07430__A1 (.DIODE(\B_type_imm[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07041__A (.DIODE(\B_type_imm[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10224__A0 (.DIODE(\B_type_imm[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07396__A (.DIODE(\B_type_imm[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07102__B1 (.DIODE(\B_type_imm[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07099__B (.DIODE(\B_type_imm[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07096__B (.DIODE(\B_type_imm[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10262__A0 (.DIODE(\B_type_imm[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07101__A (.DIODE(\B_type_imm[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07098__B (.DIODE(\B_type_imm[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10221__A0 (.DIODE(\B_type_imm[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07393__A (.DIODE(\B_type_imm[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07104__B (.DIODE(\B_type_imm[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07081__B (.DIODE(\B_type_imm[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07080__B (.DIODE(\B_type_imm[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10298__A0 (.DIODE(\B_type_imm[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07423__A (.DIODE(\B_type_imm[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07078__B (.DIODE(\B_type_imm[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07077__B (.DIODE(\B_type_imm[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07334__B (.DIODE(\J_type_imm[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07332__A (.DIODE(\J_type_imm[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07328__B (.DIODE(\J_type_imm[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07323__B_N (.DIODE(\J_type_imm[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07321__B (.DIODE(\J_type_imm[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07069__B (.DIODE(\J_type_imm[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07065__B (.DIODE(\J_type_imm[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10881__A (.DIODE(\J_type_imm[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07486__B (.DIODE(\J_type_imm[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07334__A (.DIODE(\J_type_imm[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07333__B (.DIODE(\J_type_imm[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07328__A (.DIODE(\J_type_imm[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07323__A (.DIODE(\J_type_imm[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07195__A (.DIODE(\J_type_imm[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07127__B (.DIODE(\J_type_imm[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07066__B (.DIODE(\J_type_imm[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10509__S (.DIODE(\J_type_imm[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10508__S (.DIODE(\J_type_imm[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10488__S (.DIODE(\J_type_imm[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10477__S (.DIODE(\J_type_imm[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10442__A (.DIODE(\J_type_imm[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07191__A (.DIODE(\J_type_imm[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07119__B (.DIODE(\J_type_imm[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07118__B (.DIODE(\J_type_imm[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11188__A1 (.DIODE(\J_type_imm[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07850__A0 (.DIODE(\J_type_imm[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07126__B (.DIODE(\J_type_imm[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07123__B (.DIODE(\J_type_imm[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07122__B (.DIODE(\J_type_imm[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11224__A1 (.DIODE(\J_type_imm[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07844__A0 (.DIODE(\J_type_imm[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07062__B (.DIODE(\J_type_imm[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07061__B (.DIODE(\J_type_imm[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11241__A1 (.DIODE(\J_type_imm[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07839__A0 (.DIODE(\J_type_imm[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07059__B (.DIODE(\J_type_imm[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07058__B (.DIODE(\J_type_imm[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11265__A1 (.DIODE(\J_type_imm[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07834__A0 (.DIODE(\J_type_imm[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07056__B (.DIODE(\J_type_imm[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07055__B (.DIODE(\J_type_imm[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11296__A1 (.DIODE(\J_type_imm[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07830__A1 (.DIODE(\J_type_imm[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07135__B (.DIODE(\J_type_imm[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07054__B (.DIODE(\J_type_imm[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11010__A1 (.DIODE(\PC[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09815__A0 (.DIODE(\PC[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07670__A0 (.DIODE(\PC[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07658__B1 (.DIODE(\PC[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07349__A (.DIODE(\PC[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07109__A (.DIODE(\PC[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07107__A (.DIODE(\PC[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09860__B1 (.DIODE(\PC[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07553__B2 (.DIODE(\PC[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07540__A (.DIODE(\PC[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07527__A1 (.DIODE(\PC[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07355__B (.DIODE(\PC[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07185__A1 (.DIODE(\PC[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07146__A (.DIODE(\PC[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07056__A (.DIODE(\PC[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07055__A (.DIODE(\PC[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09866__A0 (.DIODE(\PC[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07539__A2 (.DIODE(\PC[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07527__B1 (.DIODE(\PC[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07355__A (.DIODE(\PC[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07183__A (.DIODE(\PC[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07182__A (.DIODE(\PC[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07135__A (.DIODE(\PC[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07054__A (.DIODE(\PC[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11386__A1 (.DIODE(\PC[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11358__A (.DIODE(\PC[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11357__A (.DIODE(\PC[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09877__A0 (.DIODE(\PC[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07507__A2 (.DIODE(\PC[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07503__A (.DIODE(\PC[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07480__A1 (.DIODE(\PC[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07357__B (.DIODE(\PC[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07050__A (.DIODE(\PC[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07049__A (.DIODE(\PC[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11384__A (.DIODE(\PC[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11383__A (.DIODE(\PC[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09882__A0 (.DIODE(\PC[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07491__A2 (.DIODE(\PC[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07480__B1 (.DIODE(\PC[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07357__A (.DIODE(\PC[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07141__A (.DIODE(\PC[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07048__A (.DIODE(\PC[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11462__A (.DIODE(\PC[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11414__A (.DIODE(\PC[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11413__A (.DIODE(\PC[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09887__A0 (.DIODE(\PC[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07468__A1 (.DIODE(\PC[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07358__A (.DIODE(\PC[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07047__A (.DIODE(\PC[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10867__A (.DIODE(\PC[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09800__A1 (.DIODE(\PC[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07713__A2 (.DIODE(\PC[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07704__B1 (.DIODE(\PC[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07347__A (.DIODE(\PC[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07104__A (.DIODE(\PC[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07081__A (.DIODE(\PC[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07080__A (.DIODE(\PC[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10944__A1 (.DIODE(\PC[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09804__A0 (.DIODE(\PC[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07701__A0 (.DIODE(\PC[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07682__A (.DIODE(\PC[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07348__A (.DIODE(\PC[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07078__A (.DIODE(\PC[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07077__A (.DIODE(\PC[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10980__A1 (.DIODE(\PC[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09810__A0 (.DIODE(\PC[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07681__A2 (.DIODE(\PC[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07672__A (.DIODE(\PC[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07658__A1 (.DIODE(\PC[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07349__B (.DIODE(\PC[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07074__A (.DIODE(\PC[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07072__A (.DIODE(\PC[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14349__D (.DIODE(_00000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08888__B (.DIODE(_00000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08887__B (.DIODE(_00000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08885__A2 (.DIODE(_00000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08884__A1_N (.DIODE(_00000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08883__C (.DIODE(_00000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08881__A1 (.DIODE(_00000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08876__B (.DIODE(_00000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08724__B (.DIODE(_00000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14350__D (.DIODE(_00001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09697__A1 (.DIODE(_00001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09380__A1 (.DIODE(_00001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09116__A1 (.DIODE(_00001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09039__A1 (.DIODE(_00001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08717__A2 (.DIODE(_00001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08581__A1 (.DIODE(_00001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08444__A1 (.DIODE(_00001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07830__A2 (.DIODE(_00001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07803__A2 (.DIODE(_00001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14349__SET_B (.DIODE(_00068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12782__A (.DIODE(_00068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12780__A (.DIODE(_00068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12778__A (.DIODE(_00068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12776__A (.DIODE(_00068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12774__A (.DIODE(_00068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12772__A (.DIODE(_00068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12770__A (.DIODE(_00068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12768__A (.DIODE(_00068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12766__A (.DIODE(_00068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15124__D (.DIODE(_01314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15137__D (.DIODE(_01327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15220__D (.DIODE(_01410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15221__D (.DIODE(_01411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11652__C1 (.DIODE(_01527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11604__C1 (.DIODE(_01527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11559__C1 (.DIODE(_01527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11547__C1 (.DIODE(_01527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11485__C1 (.DIODE(_01527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11265__C1 (.DIODE(_01527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11010__C1 (.DIODE(_01527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10560__A (.DIODE(_01527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09740__A (.DIODE(_01527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07034__A (.DIODE(_01527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11631__C1 (.DIODE(_01528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11524__C1 (.DIODE(_01528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11440__A1 (.DIODE(_01528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11409__A1 (.DIODE(_01528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11350__A1 (.DIODE(_01528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11227__C1 (.DIODE(_01528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11049__C1 (.DIODE(_01528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10766__A (.DIODE(_01528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07628__C1 (.DIODE(_01528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07035__A (.DIODE(_01528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09731__A (.DIODE(_01529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07766__C1 (.DIODE(_01529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07618__B2 (.DIODE(_01529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07605__B1 (.DIODE(_01529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07526__A1 (.DIODE(_01529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07525__C1 (.DIODE(_01529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07491__A1 (.DIODE(_01529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07490__B1 (.DIODE(_01529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07468__A2 (.DIODE(_01529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07467__B1 (.DIODE(_01529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07463__A (.DIODE(_01531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07364__D (.DIODE(_01531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07361__A (.DIODE(_01531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07038__D (.DIODE(_01531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11011__A1 (.DIODE(_01532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10943__A1 (.DIODE(_01532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10646__A0 (.DIODE(_01532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10189__A (.DIODE(_01532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07509__B (.DIODE(_01532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07499__C1 (.DIODE(_01532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07464__A (.DIODE(_01532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07039__B (.DIODE(_01532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09725__A2 (.DIODE(_01534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07765__A (.DIODE(_01534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07680__B2 (.DIODE(_01534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07654__B1 (.DIODE(_01534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07628__A1 (.DIODE(_01534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07565__A2 (.DIODE(_01534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07544__B1 (.DIODE(_01534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07538__A2 (.DIODE(_01534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07473__B1 (.DIODE(_01534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07466__A1 (.DIODE(_01534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10435__A (.DIODE(_01535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07443__A (.DIODE(_01535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07440__A (.DIODE(_01535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07431__A1 (.DIODE(_01535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07382__A (.DIODE(_01535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07169__B (.DIODE(_01535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07168__B (.DIODE(_01535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07167__A2 (.DIODE(_01535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07166__A2 (.DIODE(_01535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07042__A (.DIODE(_01535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11653__B1 (.DIODE(_01539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11652__A1 (.DIODE(_01539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09880__A1_N (.DIODE(_01539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07635__B (.DIODE(_01539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07533__B1 (.DIODE(_01539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07469__A (.DIODE(_01539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07458__A1_N (.DIODE(_01539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07368__A (.DIODE(_01539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07141__B (.DIODE(_01539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07046__A (.DIODE(_01539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09864__A1 (.DIODE(_01540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09835__A1 (.DIODE(_01540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07785__A0 (.DIODE(_01540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07592__A1 (.DIODE(_01540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07571__A2 (.DIODE(_01540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07547__B (.DIODE(_01540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07535__A1 (.DIODE(_01540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07461__A (.DIODE(_01540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07459__A (.DIODE(_01540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07047__B (.DIODE(_01540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11386__B2 (.DIODE(_01546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11360__A1 (.DIODE(_01546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11324__A (.DIODE(_01546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09871__A (.DIODE(_01546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07526__A2 (.DIODE(_01546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07508__A (.DIODE(_01546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07356__A (.DIODE(_01546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07138__A (.DIODE(_01546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07053__A (.DIODE(_01546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11386__B1 (.DIODE(_01564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11360__A2 (.DIODE(_01564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11329__A1 (.DIODE(_01564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10615__A1 (.DIODE(_01564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10537__A (.DIODE(_01564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10215__C (.DIODE(_01564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10198__A (.DIODE(_01564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09747__A (.DIODE(_01564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07824__A0 (.DIODE(_01564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07071__B (.DIODE(_01564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12041__A2 (.DIODE(_01642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11904__B (.DIODE(_01642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11765__A_N (.DIODE(_01642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11664__B (.DIODE(_01642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10581__A (.DIODE(_01642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10576__A2 (.DIODE(_01642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09745__A (.DIODE(_01642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09744__A (.DIODE(_01642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07872__A0 (.DIODE(_01642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07149__B (.DIODE(_01642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12117__A (.DIODE(_01648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12041__A1 (.DIODE(_01648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11904__A (.DIODE(_01648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11765__C (.DIODE(_01648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11664__A (.DIODE(_01648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10582__A (.DIODE(_01648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10576__A1 (.DIODE(_01648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09720__A (.DIODE(_01648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07870__A0 (.DIODE(_01648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07155__A (.DIODE(_01648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07728__B (.DIODE(_01654_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07716__A2 (.DIODE(_01654_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07684__B (.DIODE(_01654_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07162__A4 (.DIODE(_01654_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11116__B2 (.DIODE(_01687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10802__A1 (.DIODE(_01687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10627__A (.DIODE(_01687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10608__A (.DIODE(_01687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07852__A (.DIODE(_01687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07335__A (.DIODE(_01687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07333__A (.DIODE(_01687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07330__A (.DIODE(_01687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07326__A (.DIODE(_01687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07194__A (.DIODE(_01687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11229__A1 (.DIODE(_01688_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11108__A (.DIODE(_01688_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10540__S1 (.DIODE(_01688_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10436__A (.DIODE(_01688_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10219__A (.DIODE(_01688_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07486__A (.DIODE(_01688_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07338__A (.DIODE(_01688_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07321__A (.DIODE(_01688_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07196__A (.DIODE(_01688_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11648__A1 (.DIODE(_01689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11121__A1 (.DIODE(_01689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10627__B (.DIODE(_01689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10554__A1 (.DIODE(_01689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09951__B (.DIODE(_01689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09893__A1 (.DIODE(_01689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07857__A0 (.DIODE(_01689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07475__A (.DIODE(_01689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07322__A (.DIODE(_01689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07196__B (.DIODE(_01689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07689__C1 (.DIODE(_01690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07663__C1 (.DIODE(_01690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07611__A1 (.DIODE(_01690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07598__A1 (.DIODE(_01690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07590__A1 (.DIODE(_01690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07551__A1 (.DIODE(_01690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07341__A (.DIODE(_01690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09984__A (.DIODE(_01707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09115__A (.DIODE(_01707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07214__B1 (.DIODE(_01707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10496__A0 (.DIODE(_01711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10351__A (.DIODE(_01711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10350__A (.DIODE(_01711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07240__A (.DIODE(_01711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07219__A1 (.DIODE(_01711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10516__A0 (.DIODE(_01714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10373__A (.DIODE(_01714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10372__A (.DIODE(_01714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07235__A (.DIODE(_01714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07222__A1 (.DIODE(_01714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11307__A (.DIODE(_01717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11306__A (.DIODE(_01717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10487__A0 (.DIODE(_01717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10470__A1 (.DIODE(_01717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10326__A (.DIODE(_01717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08282__A1 (.DIODE(_01717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07453__B (.DIODE(_01717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07375__A (.DIODE(_01717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07308__A1 (.DIODE(_01717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07233__A1 (.DIODE(_01717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11250__A (.DIODE(_01723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11249__A (.DIODE(_01723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10508__A0 (.DIODE(_01723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10443__A1 (.DIODE(_01723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10333__A (.DIODE(_01723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08329__A1 (.DIODE(_01723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07533__A1 (.DIODE(_01723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07450__B (.DIODE(_01723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07375__C (.DIODE(_01723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07230__B (.DIODE(_01723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11594__A (.DIODE(_01736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11562__A (.DIODE(_01736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11560__A (.DIODE(_01736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10569__B (.DIODE(_01736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10488__A1 (.DIODE(_01736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10469__A0 (.DIODE(_01736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10407__B (.DIODE(_01736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10406__A (.DIODE(_01736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08059__A0 (.DIODE(_01736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07243__A1 (.DIODE(_01736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11150__A1 (.DIODE(_01747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11100__A1 (.DIODE(_01747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10487__A1 (.DIODE(_01747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10470__A0 (.DIODE(_01747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10313__A1 (.DIODE(_01747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08443__A (.DIODE(_01747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07435__B (.DIODE(_01747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07434__B (.DIODE(_01747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07379__B (.DIODE(_01747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07264__A1 (.DIODE(_01747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11040__A (.DIODE(_01749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11039__A (.DIODE(_01749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10567__A (.DIODE(_01749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10491__A0 (.DIODE(_01749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10472__A1 (.DIODE(_01749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08466__A1 (.DIODE(_01749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07431__A2 (.DIODE(_01749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07430__A2 (.DIODE(_01749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07382__B (.DIODE(_01749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07264__B2 (.DIODE(_01749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10973__A (.DIODE(_01752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10972__A (.DIODE(_01752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10567__C (.DIODE(_01752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10512__A0 (.DIODE(_01752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10448__A1 (.DIODE(_01752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10302__A (.DIODE(_01752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08511__A1 (.DIODE(_01752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07390__B (.DIODE(_01752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07389__B (.DIODE(_01752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07259__B2 (.DIODE(_01752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11003__B2 (.DIODE(_01754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10955__A1 (.DIODE(_01754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10496__A1 (.DIODE(_01754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10309__A1 (.DIODE(_01754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07296__A (.DIODE(_01754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07261__A2_N (.DIODE(_01754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10565__D (.DIODE(_01764_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10490__A1 (.DIODE(_01764_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10473__A0 (.DIODE(_01764_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10255__A (.DIODE(_01764_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09779__B (.DIODE(_01764_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09778__B (.DIODE(_01764_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08628__A1 (.DIODE(_01764_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07401__B (.DIODE(_01764_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07399__B (.DIODE(_01764_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07271__A (.DIODE(_01764_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10892__A (.DIODE(_01767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10267__A (.DIODE(_01767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10263__A (.DIODE(_01767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08580__A (.DIODE(_01767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07274__B2 (.DIODE(_01767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10461__A (.DIODE(_01770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10451__A0 (.DIODE(_01770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09987__B2 (.DIODE(_01770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09961__B2 (.DIODE(_01770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09935__B2 (.DIODE(_01770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09916__A (.DIODE(_01770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09651__A0 (.DIODE(_01770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07316__B1 (.DIODE(_01770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07289__B1 (.DIODE(_01770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07280__A2 (.DIODE(_01770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10728__A1 (.DIODE(_01772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10466__A0 (.DIODE(_01772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09985__B2 (.DIODE(_01772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09958__B2 (.DIODE(_01772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09932__B2 (.DIODE(_01772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09914__A (.DIODE(_01772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09674__A1 (.DIODE(_01772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07317__B1 (.DIODE(_01772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07287__A2 (.DIODE(_01772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07280__B1 (.DIODE(_01772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10666__B1 (.DIODE(_01778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10564__C (.DIODE(_01778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10509__A0 (.DIODE(_01778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10441__A1 (.DIODE(_01778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10234__B1 (.DIODE(_01778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08694__A1 (.DIODE(_01778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07411__B (.DIODE(_01778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07410__B (.DIODE(_01778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07314__A1 (.DIODE(_01778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07286__A (.DIODE(_01778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09696__A (.DIODE(_01779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07314__A2 (.DIODE(_01779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07286__B (.DIODE(_01779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10884__A (.DIODE(_01784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10883__A (.DIODE(_01784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10565__A (.DIODE(_01784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10497__A0 (.DIODE(_01784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10479__A1 (.DIODE(_01784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08557__A1 (.DIODE(_01784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07427__B (.DIODE(_01784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07394__B (.DIODE(_01784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07301__A1 (.DIODE(_01784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07294__A1 (.DIODE(_01784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07318__A (.DIODE(_01794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07301__C1 (.DIODE(_01794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07319__A (.DIODE(_01803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07310__B1 (.DIODE(_01803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10667__A1 (.DIODE(_01807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10604__A (.DIODE(_01807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10564__D (.DIODE(_01807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10500__A1 (.DIODE(_01807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10238__A (.DIODE(_01807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10237__A (.DIODE(_01807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09747__B (.DIODE(_01807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09745__B (.DIODE(_01807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09744__B (.DIODE(_01807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07314__B2 (.DIODE(_01807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07339__A (.DIODE(_01813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07331__A (.DIODE(_01813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07325__B (.DIODE(_01813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07320__B1 (.DIODE(_01813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07336__A1_N (.DIODE(_01814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07327__A1 (.DIODE(_01814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11280__C1 (.DIODE(_01816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11074__A1 (.DIODE(_01816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10837__B2 (.DIODE(_01816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10805__B2 (.DIODE(_01816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10711__B1 (.DIODE(_01816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10629__A1 (.DIODE(_01816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07478__A (.DIODE(_01816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07327__A2 (.DIODE(_01816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11589__A1 (.DIODE(_01823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11540__A1 (.DIODE(_01823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11108__B (.DIODE(_01823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10863__A (.DIODE(_01823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10802__B1 (.DIODE(_01823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10747__A (.DIODE(_01823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07330__B (.DIODE(_01823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11061__A1 (.DIODE(_01826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10627__C (.DIODE(_01826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10433__A1 (.DIODE(_01826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10428__A (.DIODE(_01826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09903__A (.DIODE(_01826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09893__A2 (.DIODE(_01826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09890__A (.DIODE(_01826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07860__A0 (.DIODE(_01826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07475__B_N (.DIODE(_01826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07333__C (.DIODE(_01826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11279__A (.DIODE(_01827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11251__A1 (.DIODE(_01827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10805__A1_N (.DIODE(_01827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10712__A (.DIODE(_01827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10542__A (.DIODE(_01827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07336__A2_N (.DIODE(_01827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10651__A (.DIODE(_01828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10552__A (.DIODE(_01828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10219__B (.DIODE(_01828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07335__B (.DIODE(_01828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11466__A0 (.DIODE(_01829_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11280__A1 (.DIODE(_01829_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11145__A0 (.DIODE(_01829_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11073__A0 (.DIODE(_01829_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10925__A0 (.DIODE(_01829_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10836__A0 (.DIODE(_01829_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10711__A1 (.DIODE(_01829_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10628__A0 (.DIODE(_01829_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10541__A (.DIODE(_01829_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07336__B1 (.DIODE(_01829_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09906__A (.DIODE(_01832_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09895__A1 (.DIODE(_01832_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07607__A1 (.DIODE(_01832_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07569__A1 (.DIODE(_01832_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07339__B (.DIODE(_01832_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07688__A (.DIODE(_01836_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07662__A (.DIODE(_01836_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07637__B2 (.DIODE(_01836_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07549__B1 (.DIODE(_01836_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07517__A (.DIODE(_01836_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07516__B1 (.DIODE(_01836_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07500__A (.DIODE(_01836_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07343__A (.DIODE(_01836_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07678__S (.DIODE(_01837_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07648__S (.DIODE(_01837_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07610__A1 (.DIODE(_01837_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07586__B1 (.DIODE(_01837_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07569__B1 (.DIODE(_01837_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07557__A (.DIODE(_01837_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07531__A (.DIODE(_01837_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07485__A1 (.DIODE(_01837_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07363__B2 (.DIODE(_01837_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07344__B1 (.DIODE(_01837_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11435__A2_N (.DIODE(_01852_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07467__A1 (.DIODE(_01852_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07363__B1 (.DIODE(_01852_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10558__C (.DIODE(_01854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10269__A1 (.DIODE(_01854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10268__A (.DIODE(_01854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10231__A1 (.DIODE(_01854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10227__A1 (.DIODE(_01854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10185__D (.DIODE(_01854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10180__B (.DIODE(_01854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09734__B (.DIODE(_01854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07463__B (.DIODE(_01854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07361__B (.DIODE(_01854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07679__A (.DIODE(_01856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07649__A (.DIODE(_01856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07617__A1 (.DIODE(_01856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07590__C1 (.DIODE(_01856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07574__A (.DIODE(_01856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07559__A (.DIODE(_01856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07551__C1 (.DIODE(_01856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07524__A1 (.DIODE(_01856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07488__B1 (.DIODE(_01856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07363__C1 (.DIODE(_01856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11135__A (.DIODE(_01858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10850__A1_N (.DIODE(_01858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10811__A1_N (.DIODE(_01858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10721__A1_N (.DIODE(_01858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07365__A (.DIODE(_01858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11435__A1_N (.DIODE(_01859_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11362__A (.DIODE(_01859_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11297__A1 (.DIODE(_01859_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11255__A1 (.DIODE(_01859_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11225__A (.DIODE(_01859_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11123__A (.DIODE(_01859_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11062__A (.DIODE(_01859_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11047__A (.DIODE(_01859_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10764__A (.DIODE(_01859_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07366__A (.DIODE(_01859_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09725__B2 (.DIODE(_01861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07766__A1 (.DIODE(_01861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07699__B1 (.DIODE(_01861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07680__A1 (.DIODE(_01861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07668__A1 (.DIODE(_01861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07621__A (.DIODE(_01861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07552__A1 (.DIODE(_01861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07537__B2 (.DIODE(_01861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07489__A1 (.DIODE(_01861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07465__A1 (.DIODE(_01861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10521__A1 (.DIODE(_01867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10455__A0 (.DIODE(_01867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10369__A (.DIODE(_01867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10324__A (.DIODE(_01867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10323__A (.DIODE(_01867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09864__A2 (.DIODE(_01867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08306__A1 (.DIODE(_01867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07535__A2 (.DIODE(_01867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07452__B (.DIODE(_01867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07375__B (.DIODE(_01867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11245__A1 (.DIODE(_01868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10501__A1 (.DIODE(_01868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10476__A0 (.DIODE(_01868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10367__A1 (.DIODE(_01868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10342__A (.DIODE(_01868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08353__A1 (.DIODE(_01868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07533__A2 (.DIODE(_01868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07447__B (.DIODE(_01868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07446__B (.DIODE(_01868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07375__D (.DIODE(_01868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11199__A (.DIODE(_01870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11178__A1 (.DIODE(_01870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11177__A (.DIODE(_01870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10501__A0 (.DIODE(_01870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10476__A1 (.DIODE(_01870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10318__A (.DIODE(_01870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10314__B (.DIODE(_01870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08376__A0 (.DIODE(_01870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07443__B (.DIODE(_01870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07380__A (.DIODE(_01870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11207__A1 (.DIODE(_01871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11168__A1 (.DIODE(_01871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10508__A1 (.DIODE(_01871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10443__A0 (.DIODE(_01871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10319__A1 (.DIODE(_01871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10275__B1 (.DIODE(_01871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08399__A1 (.DIODE(_01871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07441__B (.DIODE(_01871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07440__B (.DIODE(_01871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07380__B (.DIODE(_01871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11197__A1 (.DIODE(_01872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11111__A (.DIODE(_01872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11103__A (.DIODE(_01872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10521__A0 (.DIODE(_01872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10455__A1 (.DIODE(_01872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10312__B (.DIODE(_01872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10280__B_N (.DIODE(_01872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08421__A1 (.DIODE(_01872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07438__B (.DIODE(_01872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07379__A (.DIODE(_01872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11083__A1 (.DIODE(_01877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11020__A1 (.DIODE(_01877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10567__B (.DIODE(_01877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10459__A0 (.DIODE(_01877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10310__A (.DIODE(_01877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10291__A (.DIODE(_01877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08489__A1 (.DIODE(_01877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07429__A2 (.DIODE(_01877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07386__A (.DIODE(_01877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07384__B (.DIODE(_01877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09818__B1 (.DIODE(_01881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07651__B1 (.DIODE(_01881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07430__C1 (.DIODE(_01881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07388__B (.DIODE(_01881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11601__A2 (.DIODE(_01887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11599__C (.DIODE(_01887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11547__A1 (.DIODE(_01887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11544__A (.DIODE(_01887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11543__A (.DIODE(_01887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10205__D_N (.DIODE(_01887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10199__A (.DIODE(_01887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07793__A0 (.DIODE(_01887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07427__A (.DIODE(_01887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07394__A (.DIODE(_01887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11471__A1 (.DIODE(_01892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11465__A1 (.DIODE(_01892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11463__C1 (.DIODE(_01892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10214__C (.DIODE(_01892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10205__C (.DIODE(_01892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10200__A (.DIODE(_01892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07803__A1 (.DIODE(_01892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07747__B (.DIODE(_01892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07401__A (.DIODE(_01892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07399__A (.DIODE(_01892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11462__B (.DIODE(_01897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11435__B2 (.DIODE(_01897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11414__B (.DIODE(_01897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11413__B (.DIODE(_01897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10462__A (.DIODE(_01897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10451__A1 (.DIODE(_01897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10196__A (.DIODE(_01897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07807__A0 (.DIODE(_01897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07414__A (.DIODE(_01897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07405__A (.DIODE(_01897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10730__A (.DIODE(_01898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10564__A (.DIODE(_01898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10488__A0 (.DIODE(_01898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10469__A1 (.DIODE(_01898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10241__B1 (.DIODE(_01898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09770__B (.DIODE(_01898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09769__B (.DIODE(_01898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08650__A1 (.DIODE(_01898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07414__B (.DIODE(_01898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07405__B (.DIODE(_01898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11392__A1 (.DIODE(_01900_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11384__B (.DIODE(_01900_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11383__B (.DIODE(_01900_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10728__A0 (.DIODE(_01900_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10466__A1 (.DIODE(_01900_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10214__D (.DIODE(_01900_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10197__C (.DIODE(_01900_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07812__A0 (.DIODE(_01900_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07413__A (.DIODE(_01900_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07408__A (.DIODE(_01900_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10729__A1 (.DIODE(_01901_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10564__B (.DIODE(_01901_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10520__A1 (.DIODE(_01901_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10456__A0 (.DIODE(_01901_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10251__A1 (.DIODE(_01901_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09762__B (.DIODE(_01901_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09761__B (.DIODE(_01901_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08672__A1 (.DIODE(_01901_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07413__B (.DIODE(_01901_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07408__B (.DIODE(_01901_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07700__A1 (.DIODE(_01958_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07669__A1 (.DIODE(_01958_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07605__A1 (.DIODE(_01958_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07599__B1 (.DIODE(_01958_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07525__A1 (.DIODE(_01958_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07490__A1 (.DIODE(_01958_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07489__D1 (.DIODE(_01958_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07467__A2 (.DIODE(_01958_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07465__B1 (.DIODE(_01958_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11030__C1 (.DIODE(_01970_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10991__C1 (.DIODE(_01970_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10964__C1 (.DIODE(_01970_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10873__C1 (.DIODE(_01970_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10793__C1 (.DIODE(_01970_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10754__C1 (.DIODE(_01970_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10710__C1 (.DIODE(_01970_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10619__A (.DIODE(_01970_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10554__B1 (.DIODE(_01970_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07482__A1 (.DIODE(_01970_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11563__A1 (.DIODE(_01971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11467__A1 (.DIODE(_01971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11146__A1 (.DIODE(_01971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11110__A1 (.DIODE(_01971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10999__A1 (.DIODE(_01971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10926__A1 (.DIODE(_01971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10757__A1 (.DIODE(_01971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10650__B2 (.DIODE(_01971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10543__C1 (.DIODE(_01971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07479__A (.DIODE(_01971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11623__A1 (.DIODE(_01972_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11588__B2 (.DIODE(_01972_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11516__A1 (.DIODE(_01972_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11395__A1 (.DIODE(_01972_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11319__A1 (.DIODE(_01972_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11218__A1 (.DIODE(_01972_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07607__A2 (.DIODE(_01972_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07586__A1 (.DIODE(_01972_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07516__A1 (.DIODE(_01972_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07482__A2 (.DIODE(_01972_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11393__A2 (.DIODE(_01974_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07490__A2 (.DIODE(_01974_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07487__B1 (.DIODE(_01974_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07483__B1 (.DIODE(_01974_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07482__B1 (.DIODE(_01974_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10434__A (.DIODE(_01979_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09903__B (.DIODE(_01979_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09890__B (.DIODE(_01979_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07690__A1 (.DIODE(_01979_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07664__A1 (.DIODE(_01979_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07637__C1 (.DIODE(_01979_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07606__A1 (.DIODE(_01979_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07589__C1 (.DIODE(_01979_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07546__A (.DIODE(_01979_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07487__A2 (.DIODE(_01979_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11607__B1 (.DIODE(_01984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11550__B1 (.DIODE(_01984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11408__B1 (.DIODE(_01984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11190__D1 (.DIODE(_01984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11165__B1 (.DIODE(_01984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07775__C1 (.DIODE(_01984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07600__C1 (.DIODE(_01984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07564__B1 (.DIODE(_01984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07505__A (.DIODE(_01984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07493__A (.DIODE(_01984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09727__A (.DIODE(_01985_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07750__C1 (.DIODE(_01985_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07737__C1 (.DIODE(_01985_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07725__C1 (.DIODE(_01985_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07712__C1 (.DIODE(_01985_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07701__S (.DIODE(_01985_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07670__S (.DIODE(_01985_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07655__C1 (.DIODE(_01985_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07642__S (.DIODE(_01985_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07494__A (.DIODE(_01985_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07778__A1 (.DIODE(_01986_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07767__B2 (.DIODE(_01986_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07738__A1 (.DIODE(_01986_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07713__A1 (.DIODE(_01986_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07631__B2 (.DIODE(_01986_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07602__B1 (.DIODE(_01986_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07583__B2 (.DIODE(_01986_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07566__B2 (.DIODE(_01986_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07553__B1 (.DIODE(_01986_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07507__A1 (.DIODE(_01986_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09878__A0 (.DIODE(_01988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07499__A2 (.DIODE(_01988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07776__A2 (.DIODE(_01993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07758__A (.DIODE(_01993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07751__A1 (.DIODE(_01993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07737__A1 (.DIODE(_01993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07726__A1 (.DIODE(_01993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07703__B1 (.DIODE(_01993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07506__B2 (.DIODE(_01993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07502__B (.DIODE(_01993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09727__B (.DIODE(_01994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07777__A2 (.DIODE(_01994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07754__A (.DIODE(_01994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07741__A (.DIODE(_01994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07736__A1 (.DIODE(_01994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07715__A (.DIODE(_01994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07711__A1 (.DIODE(_01994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07627__A (.DIODE(_01994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07529__A1 (.DIODE(_01994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07506__A1 (.DIODE(_01994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11362__B (.DIODE(_01995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07506__A2 (.DIODE(_01995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07752__A1 (.DIODE(_01997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07727__A1 (.DIODE(_01997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07681__A1 (.DIODE(_01997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07673__B1 (.DIODE(_01997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07657__A1 (.DIODE(_01997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07577__C1 (.DIODE(_01997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07541__B1 (.DIODE(_01997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07539__A1 (.DIODE(_01997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07529__B1 (.DIODE(_01997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07506__C1 (.DIODE(_01997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07775__B2 (.DIODE(_02000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07750__B2 (.DIODE(_02000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07735__B (.DIODE(_02000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07725__B2 (.DIODE(_02000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07710__A (.DIODE(_02000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07641__B2 (.DIODE(_02000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07615__B1 (.DIODE(_02000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07600__A1 (.DIODE(_02000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07581__B1 (.DIODE(_02000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07512__A (.DIODE(_02000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07750__A1 (.DIODE(_02013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07736__B2 (.DIODE(_02013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07725__A1 (.DIODE(_02013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07711__B2 (.DIODE(_02013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07656__A1 (.DIODE(_02013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07616__A1 (.DIODE(_02013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07601__A1 (.DIODE(_02013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07577__B2 (.DIODE(_02013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07562__A (.DIODE(_02013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07524__B2 (.DIODE(_02013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07673__A1 (.DIODE(_02014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07655__A1 (.DIODE(_02014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07617__C1 (.DIODE(_02014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07577__A1 (.DIODE(_02014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07564__A1 (.DIODE(_02014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07541__A1 (.DIODE(_02014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07524__C1 (.DIODE(_02014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09726__A2 (.DIODE(_02021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07630__B (.DIODE(_02021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07537__A1 (.DIODE(_02021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13241__A_N (.DIODE(_02241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12968__B (.DIODE(_02241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12392__C (.DIODE(_02241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12255__B (.DIODE(_02241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11835__C_N (.DIODE(_02241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11665__C (.DIODE(_02241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10585__B (.DIODE(_02241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10575__C (.DIODE(_02241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07868__A0 (.DIODE(_02241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07769__B (.DIODE(_02241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08990__B (.DIODE(_02252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07960__B (.DIODE(_02252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07882__A (.DIODE(_02252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07859__A (.DIODE(_02252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07801__B (.DIODE(_02252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07784__A (.DIODE(_02252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07781__A (.DIODE(_02252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09651__S (.DIODE(_02253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09538__S (.DIODE(_02253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09492__S (.DIODE(_02253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09312__S (.DIODE(_02253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09190__S (.DIODE(_02253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09139__S (.DIODE(_02253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08579__A (.DIODE(_02253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07828__B (.DIODE(_02253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07806__A (.DIODE(_02253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07782__A (.DIODE(_02253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09696__B (.DIODE(_02254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09605__C1 (.DIODE(_02254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09424__C1 (.DIODE(_02254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09266__C1 (.DIODE(_02254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08944__C1 (.DIODE(_02254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08627__C1 (.DIODE(_02254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08488__C1 (.DIODE(_02254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08328__C1 (.DIODE(_02254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08135__C1 (.DIODE(_02254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07783__A (.DIODE(_02254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09070__A (.DIODE(_02255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08330__A (.DIODE(_02255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07889__A (.DIODE(_02255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07797__S (.DIODE(_02255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07795__S (.DIODE(_02255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07793__S (.DIODE(_02255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07791__S (.DIODE(_02255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07789__S (.DIODE(_02255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07787__S (.DIODE(_02255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07785__S (.DIODE(_02255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09650__A1 (.DIODE(_02263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09603__B1 (.DIODE(_02263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09537__A1 (.DIODE(_02263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09422__B1 (.DIODE(_02263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09264__B1 (.DIODE(_02263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08942__B1 (.DIODE(_02263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07800__A (.DIODE(_02263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09687__C1 (.DIODE(_02264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09491__A1 (.DIODE(_02264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09370__C1 (.DIODE(_02264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09311__A1 (.DIODE(_02264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09189__A1 (.DIODE(_02264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09138__A1 (.DIODE(_02264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09106__C1 (.DIODE(_02264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09067__A1 (.DIODE(_02264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09021__C1 (.DIODE(_02264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07801__A (.DIODE(_02264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09719__B1 (.DIODE(_02265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09674__B1 (.DIODE(_02265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09628__B1 (.DIODE(_02265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09583__B1 (.DIODE(_02265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09561__B1 (.DIODE(_02265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09515__B1 (.DIODE(_02265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09469__B1 (.DIODE(_02265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09447__B1 (.DIODE(_02265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07802__A (.DIODE(_02265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09402__B1 (.DIODE(_02266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09357__B1 (.DIODE(_02266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09335__B1 (.DIODE(_02266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09289__B1 (.DIODE(_02266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09244__B1 (.DIODE(_02266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09216__B1 (.DIODE(_02266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09167__B1 (.DIODE(_02266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09093__B1 (.DIODE(_02266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08993__B1 (.DIODE(_02266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07803__B1 (.DIODE(_02266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09645__C1 (.DIODE(_02267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09587__B1 (.DIODE(_02267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09532__C1 (.DIODE(_02267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09486__C1 (.DIODE(_02267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09406__B1 (.DIODE(_02267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09306__C1 (.DIODE(_02267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09248__B1 (.DIODE(_02267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09019__A (.DIODE(_02267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08906__B1 (.DIODE(_02267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07805__A (.DIODE(_02267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09717__A1 (.DIODE(_02268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09513__C1 (.DIODE(_02268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09355__A1 (.DIODE(_02268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09333__A1 (.DIODE(_02268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09287__A1 (.DIODE(_02268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09214__A1 (.DIODE(_02268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09164__C1 (.DIODE(_02268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09091__A1 (.DIODE(_02268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08991__A1 (.DIODE(_02268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07807__A1 (.DIODE(_02268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07857__S (.DIODE(_02269_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07855__S (.DIODE(_02269_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07850__S (.DIODE(_02269_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07844__S (.DIODE(_02269_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07839__S (.DIODE(_02269_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07834__S (.DIODE(_02269_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07824__S (.DIODE(_02269_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07818__S (.DIODE(_02269_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07812__S (.DIODE(_02269_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07807__S (.DIODE(_02269_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09644__A (.DIODE(_02271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09531__A (.DIODE(_02271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09485__A (.DIODE(_02271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09305__A (.DIODE(_02271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09183__A (.DIODE(_02271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09132__A (.DIODE(_02271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09065__S (.DIODE(_02271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09059__A (.DIODE(_02271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09017__A (.DIODE(_02271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07810__A (.DIODE(_02271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09594__S (.DIODE(_02272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09512__C1 (.DIODE(_02272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09413__S (.DIODE(_02272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09255__S (.DIODE(_02272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09163__C1 (.DIODE(_02272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09129__A1 (.DIODE(_02272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09054__A1 (.DIODE(_02272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08975__A (.DIODE(_02272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08923__S (.DIODE(_02272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07811__A (.DIODE(_02272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09659__A1 (.DIODE(_02273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09613__A1 (.DIODE(_02273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09568__A1 (.DIODE(_02273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09546__A1 (.DIODE(_02273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09454__A1 (.DIODE(_02273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09432__A1 (.DIODE(_02273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09387__A1 (.DIODE(_02273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09227__A1 (.DIODE(_02273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08957__A1 (.DIODE(_02273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07812__A1 (.DIODE(_02273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11356__A1 (.DIODE(_02276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09600__B1 (.DIODE(_02276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09419__B1 (.DIODE(_02276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09261__B1 (.DIODE(_02276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09219__A (.DIODE(_02276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09031__A (.DIODE(_02276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08937__B1 (.DIODE(_02276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08926__A (.DIODE(_02276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08920__A (.DIODE(_02276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07816__A (.DIODE(_02276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09710__B1 (.DIODE(_02277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09693__S1 (.DIODE(_02277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09376__S1 (.DIODE(_02277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09352__B1 (.DIODE(_02277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09326__B1 (.DIODE(_02277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09280__B1 (.DIODE(_02277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09205__B1 (.DIODE(_02277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09088__B1 (.DIODE(_02277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08985__B1 (.DIODE(_02277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07817__A (.DIODE(_02277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09716__A1 (.DIODE(_02278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09395__A1 (.DIODE(_02278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09350__A1 (.DIODE(_02278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09332__A1 (.DIODE(_02278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09286__A1 (.DIODE(_02278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09236__A1 (.DIODE(_02278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09213__A1 (.DIODE(_02278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09086__A1 (.DIODE(_02278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08982__A1 (.DIODE(_02278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07818__A1 (.DIODE(_02278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09639__S0 (.DIODE(_02280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09526__S0 (.DIODE(_02280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09480__S0 (.DIODE(_02280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09047__A (.DIODE(_02280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09045__A (.DIODE(_02280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09009__A (.DIODE(_02280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09002__A (.DIODE(_02280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08958__A (.DIODE(_02280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08938__A (.DIODE(_02280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07821__A (.DIODE(_02280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09635__S (.DIODE(_02281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09522__S (.DIODE(_02281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09476__S (.DIODE(_02281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09304__S0 (.DIODE(_02281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09296__S (.DIODE(_02281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09182__S0 (.DIODE(_02281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09131__S0 (.DIODE(_02281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09058__S0 (.DIODE(_02281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08919__A (.DIODE(_02281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07822__A (.DIODE(_02281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09593__S0 (.DIODE(_02282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09592__S0 (.DIODE(_02282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09412__S0 (.DIODE(_02282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09303__S0 (.DIODE(_02282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09254__S0 (.DIODE(_02282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09181__S0 (.DIODE(_02282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09130__S0 (.DIODE(_02282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09057__S0 (.DIODE(_02282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08922__S0 (.DIODE(_02282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07823__A (.DIODE(_02282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09706__S0 (.DIODE(_02283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09344__S0 (.DIODE(_02283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09322__S0 (.DIODE(_02283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09276__S0 (.DIODE(_02283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09200__S0 (.DIODE(_02283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09081__S0 (.DIODE(_02283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09079__S0 (.DIODE(_02283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08974__S0 (.DIODE(_02283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08973__S0 (.DIODE(_02283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07824__A1 (.DIODE(_02283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08706__B1 (.DIODE(_02285_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08625__B1 (.DIODE(_02285_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08486__B1 (.DIODE(_02285_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08326__B1 (.DIODE(_02285_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07827__A (.DIODE(_02285_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08603__A1 (.DIODE(_02286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08570__C1 (.DIODE(_02286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08533__A1 (.DIODE(_02286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08434__C1 (.DIODE(_02286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08375__A1 (.DIODE(_02286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08258__A1 (.DIODE(_02286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08133__B1 (.DIODE(_02286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08058__A1 (.DIODE(_02286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07997__A1 (.DIODE(_02286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07828__A (.DIODE(_02286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08282__B1 (.DIODE(_02288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08236__B1 (.DIODE(_02288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08213__B1 (.DIODE(_02288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08189__B1 (.DIODE(_02288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08167__B1 (.DIODE(_02288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08109__B1 (.DIODE(_02288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08084__B1 (.DIODE(_02288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08036__B1 (.DIODE(_02288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07963__B1 (.DIODE(_02288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07830__B1 (.DIODE(_02288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08711__B1 (.DIODE(_02289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08590__C1 (.DIODE(_02289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08520__C1 (.DIODE(_02289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08362__C1 (.DIODE(_02289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08245__C1 (.DIODE(_02289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08154__A (.DIODE(_02289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08045__C1 (.DIODE(_02289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07978__C1 (.DIODE(_02289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07907__A (.DIODE(_02289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07832__A (.DIODE(_02289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08706__A1 (.DIODE(_02290_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08692__A (.DIODE(_02290_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08625__A1 (.DIODE(_02290_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08574__B1 (.DIODE(_02290_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08486__A1 (.DIODE(_02290_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08438__B1 (.DIODE(_02290_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08326__A1 (.DIODE(_02290_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08133__A1 (.DIODE(_02290_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07989__C1 (.DIODE(_02290_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07833__A (.DIODE(_02290_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08464__A1 (.DIODE(_02291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08419__A1 (.DIODE(_02291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08397__A1 (.DIODE(_02291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08304__A1 (.DIODE(_02291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08280__A1 (.DIODE(_02291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08211__A1 (.DIODE(_02291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08107__A1 (.DIODE(_02291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08082__A1 (.DIODE(_02291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07961__A1 (.DIODE(_02291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07834__A1 (.DIODE(_02291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08705__C1 (.DIODE(_02293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08597__A (.DIODE(_02293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08527__A (.DIODE(_02293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08369__A (.DIODE(_02293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08252__A (.DIODE(_02293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08080__A (.DIODE(_02293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08052__A (.DIODE(_02293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07988__A (.DIODE(_02293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07936__A (.DIODE(_02293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07837__A (.DIODE(_02293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08609__A1 (.DIODE(_02294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08508__C1 (.DIODE(_02294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08477__S (.DIODE(_02294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08350__C1 (.DIODE(_02294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08317__S (.DIODE(_02294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08233__C1 (.DIODE(_02294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08193__A (.DIODE(_02294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08124__S (.DIODE(_02294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08030__C1 (.DIODE(_02294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07838__A (.DIODE(_02294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08679__A1 (.DIODE(_02295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08657__A1 (.DIODE(_02295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08635__A1 (.DIODE(_02295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08174__A1 (.DIODE(_02295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08148__A1 (.DIODE(_02295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08088__A1 (.DIODE(_02295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08064__A1 (.DIODE(_02295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08003__A1 (.DIODE(_02295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07908__A1 (.DIODE(_02295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07839__A1 (.DIODE(_02295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11231__A1 (.DIODE(_02297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08713__S1 (.DIODE(_02297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08712__S1 (.DIODE(_02297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08710__S1 (.DIODE(_02297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08708__S1 (.DIODE(_02297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08700__A (.DIODE(_02297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08140__A (.DIODE(_02297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08130__B1 (.DIODE(_02297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07943__A (.DIODE(_02297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07842__A (.DIODE(_02297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08620__A1 (.DIODE(_02298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08571__S1 (.DIODE(_02298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08536__S1 (.DIODE(_02298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08481__A1 (.DIODE(_02298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08435__S1 (.DIODE(_02298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08321__A1 (.DIODE(_02298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08168__S1 (.DIODE(_02298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08138__S1 (.DIODE(_02298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08128__A1 (.DIODE(_02298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07843__A (.DIODE(_02298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08463__A1 (.DIODE(_02299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08418__A1 (.DIODE(_02299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08392__A1 (.DIODE(_02299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08303__A1 (.DIODE(_02299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08275__A1 (.DIODE(_02299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08210__A1 (.DIODE(_02299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08106__A1 (.DIODE(_02299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08076__A1 (.DIODE(_02299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07959__A1 (.DIODE(_02299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07844__A1 (.DIODE(_02299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08699__S (.DIODE(_02301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08592__S0 (.DIODE(_02301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08522__S0 (.DIODE(_02301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08021__A (.DIODE(_02301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07990__A (.DIODE(_02301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07968__A (.DIODE(_02301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07965__A (.DIODE(_02301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07941__A (.DIODE(_02301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07915__A (.DIODE(_02301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07847__A (.DIODE(_02301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08588__S (.DIODE(_02302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08518__S (.DIODE(_02302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08360__S (.DIODE(_02302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08243__S (.DIODE(_02302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08120__A (.DIODE(_02302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08043__S (.DIODE(_02302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07987__S0 (.DIODE(_02302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07974__S (.DIODE(_02302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07932__A (.DIODE(_02302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07848__A (.DIODE(_02302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08615__S0 (.DIODE(_02303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08614__S0 (.DIODE(_02303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08476__S0 (.DIODE(_02303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08475__S0 (.DIODE(_02303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08316__S0 (.DIODE(_02303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08250__S0 (.DIODE(_02303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08123__S0 (.DIODE(_02303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08050__S0 (.DIODE(_02303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07986__S0 (.DIODE(_02303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07849__A (.DIODE(_02303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08453__S0 (.DIODE(_02304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08408__S0 (.DIODE(_02304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08386__S0 (.DIODE(_02304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08293__S0 (.DIODE(_02304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08269__S0 (.DIODE(_02304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08200__S0 (.DIODE(_02304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08095__S0 (.DIODE(_02304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08069__S0 (.DIODE(_02304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07931__S0 (.DIODE(_02304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07850__A1 (.DIODE(_02304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11373__A (.DIODE(_02306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11305__A (.DIODE(_02306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11281__A1 (.DIODE(_02306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11253__A1 (.DIODE(_02306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11075__B2 (.DIODE(_02306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10971__A (.DIODE(_02306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10908__A (.DIODE(_02306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10652__A (.DIODE(_02306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10630__A1 (.DIODE(_02306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07853__A (.DIODE(_02306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11649__B2 (.DIODE(_02308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11589__B1 (.DIODE(_02308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11541__B2 (.DIODE(_02308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11494__A (.DIODE(_02308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11419__A (.DIODE(_02308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11181__A1 (.DIODE(_02308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11043__A1 (.DIODE(_02308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09951__A (.DIODE(_02308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09893__D1 (.DIODE(_02308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07855__A0 (.DIODE(_02308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13241__C (.DIODE(_02313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12968__D (.DIODE(_02313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12392__A (.DIODE(_02313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12255__D_N (.DIODE(_02313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11835__B (.DIODE(_02313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11665__A_N (.DIODE(_02313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10585__A (.DIODE(_02313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10575__A (.DIODE(_02313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09779__A (.DIODE(_02313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07863__A0 (.DIODE(_02313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13241__D (.DIODE(_02315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12968__A_N (.DIODE(_02315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12392__B (.DIODE(_02315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12255__A (.DIODE(_02315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11665__B_N (.DIODE(_02315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10584__A (.DIODE(_02315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10575__B (.DIODE(_02315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09770__A (.DIODE(_02315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09769__A (.DIODE(_02315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07866__A0 (.DIODE(_02315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09068__S (.DIODE(_02324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08604__S (.DIODE(_02324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08534__S (.DIODE(_02324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08376__S (.DIODE(_02324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08259__S (.DIODE(_02324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08059__S (.DIODE(_02324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07998__S (.DIODE(_02324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07887__S (.DIODE(_02324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07885__S (.DIODE(_02324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07883__S (.DIODE(_02324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08306__A2 (.DIODE(_02328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08282__A2 (.DIODE(_02328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08236__A2 (.DIODE(_02328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08213__A2 (.DIODE(_02328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08189__A2 (.DIODE(_02328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08167__A2 (.DIODE(_02328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08109__A2 (.DIODE(_02328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08084__A2 (.DIODE(_02328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08036__A2 (.DIODE(_02328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07963__A2 (.DIODE(_02328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08709__A (.DIODE(_02330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08607__A (.DIODE(_02330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08468__A (.DIODE(_02330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08391__B1 (.DIODE(_02330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08308__A (.DIODE(_02330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08274__B1 (.DIODE(_02330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08190__A (.DIODE(_02330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08075__B1 (.DIODE(_02330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07958__B1 (.DIODE(_02330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07892__A (.DIODE(_02330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08677__A (.DIODE(_02331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08655__A (.DIODE(_02331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08633__A (.DIODE(_02331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08542__A1 (.DIODE(_02331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08172__A (.DIODE(_02331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08146__A (.DIODE(_02331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08086__A (.DIODE(_02331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08062__A (.DIODE(_02331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08001__A (.DIODE(_02331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07900__A (.DIODE(_02331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08600__S0 (.DIODE(_02332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08599__S0 (.DIODE(_02332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08530__S0 (.DIODE(_02332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08372__S0 (.DIODE(_02332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08255__S0 (.DIODE(_02332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08055__S0 (.DIODE(_02332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08008__A (.DIODE(_02332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07993__S0 (.DIODE(_02332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07901__A (.DIODE(_02332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07894__A (.DIODE(_02332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08703__A1 (.DIODE(_02333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08702__B_N (.DIODE(_02333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08622__A1 (.DIODE(_02333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08483__A1 (.DIODE(_02333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08323__A1 (.DIODE(_02333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08273__S (.DIODE(_02333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08130__A1 (.DIODE(_02333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08074__S (.DIODE(_02333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08012__A (.DIODE(_02333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07895__A (.DIODE(_02333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08394__A1 (.DIODE(_02334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08284__S0 (.DIODE(_02334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08277__A1 (.DIODE(_02334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08261__S0 (.DIODE(_02334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08215__S0 (.DIODE(_02334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08191__S0 (.DIODE(_02334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08085__S0 (.DIODE(_02334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08061__S0 (.DIODE(_02334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08000__S0 (.DIODE(_02334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07899__S0 (.DIODE(_02334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08592__S1 (.DIODE(_02335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08587__B1 (.DIODE(_02335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08522__S1 (.DIODE(_02335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08517__B1 (.DIODE(_02335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08364__S1 (.DIODE(_02335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08247__S1 (.DIODE(_02335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08047__S1 (.DIODE(_02335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07981__S1 (.DIODE(_02335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07912__A (.DIODE(_02335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07897__A (.DIODE(_02335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08611__S1 (.DIODE(_02336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08610__S1 (.DIODE(_02336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08472__S1 (.DIODE(_02336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08471__S1 (.DIODE(_02336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08312__S1 (.DIODE(_02336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08311__S1 (.DIODE(_02336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08116__S1 (.DIODE(_02336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08115__S1 (.DIODE(_02336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08017__A (.DIODE(_02336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07898__A (.DIODE(_02336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08682__S1 (.DIODE(_02337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08660__S1 (.DIODE(_02337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08638__S1 (.DIODE(_02337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08545__S1 (.DIODE(_02337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08499__S1 (.DIODE(_02337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08191__S1 (.DIODE(_02337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08085__S1 (.DIODE(_02337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08061__S1 (.DIODE(_02337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08000__S1 (.DIODE(_02337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07899__S1 (.DIODE(_02337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08610__S0 (.DIODE(_02340_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08606__S0 (.DIODE(_02340_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08471__S0 (.DIODE(_02340_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08467__S0 (.DIODE(_02340_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08311__S0 (.DIODE(_02340_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08307__S0 (.DIODE(_02340_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08115__S0 (.DIODE(_02340_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08111__S0 (.DIODE(_02340_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07939__A (.DIODE(_02340_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07902__A (.DIODE(_02340_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08678__S0 (.DIODE(_02341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08656__S0 (.DIODE(_02341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08634__S0 (.DIODE(_02341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08541__S0 (.DIODE(_02341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08194__S0 (.DIODE(_02341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08173__S0 (.DIODE(_02341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08087__S0 (.DIODE(_02341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08063__S0 (.DIODE(_02341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08002__S0 (.DIODE(_02341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07906__S0 (.DIODE(_02341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08600__S1 (.DIODE(_02342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08530__S1 (.DIODE(_02342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08372__S1 (.DIODE(_02342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08359__B1 (.DIODE(_02342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08255__S1 (.DIODE(_02342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08242__B1 (.DIODE(_02342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08055__S1 (.DIODE(_02342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08042__B1 (.DIODE(_02342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07973__B1 (.DIODE(_02342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07904__A (.DIODE(_02342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08696__S1 (.DIODE(_02343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08695__S1 (.DIODE(_02343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08606__S1 (.DIODE(_02343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08467__S1 (.DIODE(_02343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08307__S1 (.DIODE(_02343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08144__A (.DIODE(_02343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08111__S1 (.DIODE(_02343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08013__A (.DIODE(_02343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08010__A (.DIODE(_02343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07905__A (.DIODE(_02343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08678__S1 (.DIODE(_02344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08656__S1 (.DIODE(_02344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08634__S1 (.DIODE(_02344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08541__S1 (.DIODE(_02344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08173__S1 (.DIODE(_02344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08147__S1 (.DIODE(_02344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08087__S1 (.DIODE(_02344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08063__S1 (.DIODE(_02344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08002__S1 (.DIODE(_02344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07906__S1 (.DIODE(_02344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08569__C1 (.DIODE(_02346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08433__C1 (.DIODE(_02346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08287__B1 (.DIODE(_02346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08264__B1 (.DIODE(_02346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08218__B1 (.DIODE(_02346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08195__B1 (.DIODE(_02346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08088__B1 (.DIODE(_02346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08064__B1 (.DIODE(_02346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08003__B1 (.DIODE(_02346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07908__B1 (.DIODE(_02346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08618__S (.DIODE(_02348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08479__S (.DIODE(_02348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08364__S0 (.DIODE(_02348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08319__S (.DIODE(_02348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08247__S0 (.DIODE(_02348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08126__S (.DIODE(_02348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08047__S0 (.DIODE(_02348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07981__S0 (.DIODE(_02348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07956__A (.DIODE(_02348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07910__A (.DIODE(_02348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08617__S (.DIODE(_02349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08591__S0 (.DIODE(_02349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08521__S0 (.DIODE(_02349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08478__S (.DIODE(_02349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08363__S0 (.DIODE(_02349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08346__A (.DIODE(_02349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08318__S (.DIODE(_02349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08125__S (.DIODE(_02349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07953__A (.DIODE(_02349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07911__A (.DIODE(_02349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08573__S0 (.DIODE(_02350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08490__S0 (.DIODE(_02350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08445__S0 (.DIODE(_02350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08437__S0 (.DIODE(_02350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08400__S0 (.DIODE(_02350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08378__S0 (.DIODE(_02350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08331__S0 (.DIODE(_02350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08065__S0 (.DIODE(_02350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08004__S0 (.DIODE(_02350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07914__S0 (.DIODE(_02350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08591__S1 (.DIODE(_02351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08521__S1 (.DIODE(_02351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08363__S1 (.DIODE(_02351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08289__A (.DIODE(_02351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08246__S1 (.DIODE(_02351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08214__A (.DIODE(_02351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08046__S1 (.DIODE(_02351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07979__S1 (.DIODE(_02351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07917__A (.DIODE(_02351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07913__A (.DIODE(_02351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08382__S1 (.DIODE(_02352_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08335__S1 (.DIODE(_02352_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08288__S1 (.DIODE(_02352_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08265__S1 (.DIODE(_02352_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08219__S1 (.DIODE(_02352_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08196__S1 (.DIODE(_02352_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08090__S1 (.DIODE(_02352_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08065__S1 (.DIODE(_02352_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08004__S1 (.DIODE(_02352_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07914__S1 (.DIODE(_02352_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08710__S0 (.DIODE(_02354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08698__S (.DIODE(_02354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08548__S (.DIODE(_02354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08180__S (.DIODE(_02354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08157__S (.DIODE(_02354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08139__A (.DIODE(_02354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08089__A (.DIODE(_02354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08025__A (.DIODE(_02354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07945__A (.DIODE(_02354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07916__A (.DIODE(_02354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08383__S0 (.DIODE(_02355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08336__S0 (.DIODE(_02355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08290__S0 (.DIODE(_02355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08266__S0 (.DIODE(_02355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08220__S0 (.DIODE(_02355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08197__S0 (.DIODE(_02355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08091__S0 (.DIODE(_02355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08066__S0 (.DIODE(_02355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08005__S0 (.DIODE(_02355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07918__S0 (.DIODE(_02355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08494__S1 (.DIODE(_02356_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08449__S1 (.DIODE(_02356_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08404__S1 (.DIODE(_02356_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08266__S1 (.DIODE(_02356_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08220__S1 (.DIODE(_02356_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08197__S1 (.DIODE(_02356_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08091__S1 (.DIODE(_02356_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08066__S1 (.DIODE(_02356_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08005__S1 (.DIODE(_02356_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07918__S1 (.DIODE(_02356_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08714__S (.DIODE(_02358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08711__A1 (.DIODE(_02358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08624__C1 (.DIODE(_02358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08612__S (.DIODE(_02358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08485__C1 (.DIODE(_02358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08325__C1 (.DIODE(_02358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08132__C1 (.DIODE(_02358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08092__A (.DIODE(_02358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07951__A (.DIODE(_02358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07920__A (.DIODE(_02358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08683__S (.DIODE(_02359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08661__S (.DIODE(_02359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08639__S (.DIODE(_02359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08574__A1 (.DIODE(_02359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08546__S (.DIODE(_02359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08178__S (.DIODE(_02359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08153__S (.DIODE(_02359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08067__S (.DIODE(_02359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08006__S (.DIODE(_02359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07921__S (.DIODE(_02359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08602__A1 (.DIODE(_02361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08594__C1 (.DIODE(_02361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08532__A1 (.DIODE(_02361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08524__C1 (.DIODE(_02361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08366__C1 (.DIODE(_02361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08249__C1 (.DIODE(_02361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08049__C1 (.DIODE(_02361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07983__C1 (.DIODE(_02361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07926__A (.DIODE(_02361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07923__A (.DIODE(_02361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08715__B2 (.DIODE(_02362_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08613__B2 (.DIODE(_02362_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08474__B2 (.DIODE(_02362_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08374__A1 (.DIODE(_02362_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08257__A1 (.DIODE(_02362_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08150__A (.DIODE(_02362_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08137__A (.DIODE(_02362_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08057__A1 (.DIODE(_02362_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07996__A1 (.DIODE(_02362_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07924__A (.DIODE(_02362_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08570__A1 (.DIODE(_02363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08338__B2 (.DIODE(_02363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08292__B2 (.DIODE(_02363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08268__B2 (.DIODE(_02363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08222__B2 (.DIODE(_02363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08199__B2 (.DIODE(_02363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08094__B2 (.DIODE(_02363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08068__B2 (.DIODE(_02363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08007__B2 (.DIODE(_02363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07925__B2 (.DIODE(_02363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07963__B2 (.DIODE(_02364_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08707__A1 (.DIODE(_02365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08626__A1 (.DIODE(_02365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08578__B2 (.DIODE(_02365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08487__A1 (.DIODE(_02365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08442__B2 (.DIODE(_02365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08327__A1 (.DIODE(_02365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08314__B2 (.DIODE(_02365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08134__A1 (.DIODE(_02365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08119__B2 (.DIODE(_02365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07927__A (.DIODE(_02365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08465__A1 (.DIODE(_02366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08420__A1 (.DIODE(_02366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08398__A1 (.DIODE(_02366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08305__A1 (.DIODE(_02366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08281__A1 (.DIODE(_02366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08212__A1 (.DIODE(_02366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08108__A1 (.DIODE(_02366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08083__A1 (.DIODE(_02366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08035__A1 (.DIODE(_02366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07962__A1 (.DIODE(_02366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08703__B1 (.DIODE(_02367_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08622__B1 (.DIODE(_02367_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08483__B1 (.DIODE(_02367_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08323__B1 (.DIODE(_02367_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08251__S1 (.DIODE(_02367_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08122__A (.DIODE(_02367_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08051__S1 (.DIODE(_02367_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07987__S1 (.DIODE(_02367_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07985__A (.DIODE(_02367_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07929__A (.DIODE(_02367_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08506__B1 (.DIODE(_02368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08394__B1 (.DIODE(_02368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08348__B1 (.DIODE(_02368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08315__S1 (.DIODE(_02368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08277__B1 (.DIODE(_02368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08231__B1 (.DIODE(_02368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08121__S1 (.DIODE(_02368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08027__B1 (.DIODE(_02368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07934__A (.DIODE(_02368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07930__A (.DIODE(_02368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08562__A (.DIODE(_02369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08426__A (.DIODE(_02369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08408__S1 (.DIODE(_02369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08386__S1 (.DIODE(_02369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08293__S1 (.DIODE(_02369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08269__S1 (.DIODE(_02369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08200__S1 (.DIODE(_02369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08095__S1 (.DIODE(_02369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08069__S1 (.DIODE(_02369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07931__S1 (.DIODE(_02369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08696__S0 (.DIODE(_02371_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08695__S0 (.DIODE(_02371_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08608__S0 (.DIODE(_02371_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08595__S0 (.DIODE(_02371_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08525__S0 (.DIODE(_02371_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08469__S0 (.DIODE(_02371_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08367__S0 (.DIODE(_02371_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08309__S0 (.DIODE(_02371_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08113__S0 (.DIODE(_02371_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07933__A (.DIODE(_02371_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08454__S0 (.DIODE(_02372_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08409__S0 (.DIODE(_02372_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08387__S0 (.DIODE(_02372_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08294__S0 (.DIODE(_02372_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08270__S0 (.DIODE(_02372_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08201__S0 (.DIODE(_02372_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08147__S0 (.DIODE(_02372_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08096__S0 (.DIODE(_02372_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08070__S0 (.DIODE(_02372_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07935__S0 (.DIODE(_02372_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08454__S1 (.DIODE(_02373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08453__S1 (.DIODE(_02373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08409__S1 (.DIODE(_02373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08387__S1 (.DIODE(_02373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08294__S1 (.DIODE(_02373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08270__S1 (.DIODE(_02373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08201__S1 (.DIODE(_02373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08096__S1 (.DIODE(_02373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08070__S1 (.DIODE(_02373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07935__S1 (.DIODE(_02373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08697__S (.DIODE(_02375_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08616__S (.DIODE(_02375_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08594__A1 (.DIODE(_02375_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08524__A1 (.DIODE(_02375_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08432__C1 (.DIODE(_02375_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08366__A1 (.DIODE(_02375_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08249__A1 (.DIODE(_02375_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08049__A1 (.DIODE(_02375_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07983__A1 (.DIODE(_02375_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07937__A (.DIODE(_02375_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08455__S (.DIODE(_02376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08438__A1 (.DIODE(_02376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08410__S (.DIODE(_02376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08388__S (.DIODE(_02376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08295__S (.DIODE(_02376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08271__S (.DIODE(_02376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08202__S (.DIODE(_02376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08097__S (.DIODE(_02376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08071__S (.DIODE(_02376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07938__S (.DIODE(_02376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08682__S0 (.DIODE(_02378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08660__S0 (.DIODE(_02378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08638__S0 (.DIODE(_02378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08545__S0 (.DIODE(_02378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08456__B_N (.DIODE(_02378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08411__B_N (.DIODE(_02378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08296__B_N (.DIODE(_02378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08203__B_N (.DIODE(_02378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08098__B_N (.DIODE(_02378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07940__B_N (.DIODE(_02378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08586__B_N (.DIODE(_02380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08516__B_N (.DIODE(_02380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08358__B_N (.DIODE(_02380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08241__B_N (.DIODE(_02380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08160__A (.DIODE(_02380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08042__A1 (.DIODE(_02380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08041__B_N (.DIODE(_02380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07973__A1 (.DIODE(_02380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07972__B_N (.DIODE(_02380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07942__A (.DIODE(_02380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08457__A1 (.DIODE(_02381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08412__A1 (.DIODE(_02381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08393__B_N (.DIODE(_02381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08297__A1 (.DIODE(_02381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08276__B_N (.DIODE(_02381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08204__A1 (.DIODE(_02381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08099__A1 (.DIODE(_02381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08078__A1 (.DIODE(_02381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08077__B_N (.DIODE(_02381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07944__A1 (.DIODE(_02381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08576__S1 (.DIODE(_02382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08575__S1 (.DIODE(_02382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08457__B1 (.DIODE(_02382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08440__S1 (.DIODE(_02382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08412__B1 (.DIODE(_02382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08297__B1 (.DIODE(_02382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08204__B1 (.DIODE(_02382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08099__B1 (.DIODE(_02382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08078__B1 (.DIODE(_02382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07944__B1 (.DIODE(_02382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08689__A1 (.DIODE(_02384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08688__B_N (.DIODE(_02384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08667__A1 (.DIODE(_02384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08666__B_N (.DIODE(_02384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08645__A1 (.DIODE(_02384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08552__A1 (.DIODE(_02384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08184__A1 (.DIODE(_02384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08162__A1 (.DIODE(_02384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08100__S (.DIODE(_02384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07946__S (.DIODE(_02384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08619__A1 (.DIODE(_02387_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08589__B2 (.DIODE(_02387_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08519__B2 (.DIODE(_02387_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08480__A1 (.DIODE(_02387_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08320__A1 (.DIODE(_02387_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08127__A1 (.DIODE(_02387_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08073__A (.DIODE(_02387_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07975__A (.DIODE(_02387_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07955__A (.DIODE(_02387_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07949__A (.DIODE(_02387_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08705__B2 (.DIODE(_02388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08686__A1 (.DIODE(_02388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08664__A1 (.DIODE(_02388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08642__A1 (.DIODE(_02388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08624__B2 (.DIODE(_02388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08485__B2 (.DIODE(_02388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08325__B2 (.DIODE(_02388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08132__B2 (.DIODE(_02388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07971__A1 (.DIODE(_02388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07950__A (.DIODE(_02388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08504__A1 (.DIODE(_02389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08459__B2 (.DIODE(_02389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08414__B2 (.DIODE(_02389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08345__A1 (.DIODE(_02389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08299__B2 (.DIODE(_02389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08229__A1 (.DIODE(_02389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08206__B2 (.DIODE(_02389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08101__B2 (.DIODE(_02389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08024__A1 (.DIODE(_02389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07952__B2 (.DIODE(_02389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08675__S (.DIODE(_02390_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08653__S (.DIODE(_02390_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08577__S (.DIODE(_02390_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08560__S (.DIODE(_02390_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08538__S (.DIODE(_02390_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08441__S (.DIODE(_02390_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08424__S (.DIODE(_02390_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08170__S (.DIODE(_02390_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08101__C1 (.DIODE(_02390_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07952__C1 (.DIODE(_02390_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08495__S0 (.DIODE(_02392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08450__S0 (.DIODE(_02392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08405__S0 (.DIODE(_02392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08389__S (.DIODE(_02392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08300__S (.DIODE(_02392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08272__S (.DIODE(_02392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08207__S (.DIODE(_02392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08102__S (.DIODE(_02392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08072__S (.DIODE(_02392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07954__S (.DIODE(_02392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08701__A1 (.DIODE(_02394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08549__A1 (.DIODE(_02394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08462__A1 (.DIODE(_02394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08417__A1 (.DIODE(_02394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08302__A1 (.DIODE(_02394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08209__A1 (.DIODE(_02394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08181__A1 (.DIODE(_02394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08158__A1 (.DIODE(_02394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08105__A1 (.DIODE(_02394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07958__A1 (.DIODE(_02394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08461__S (.DIODE(_02395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08416__S (.DIODE(_02395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08390__S (.DIODE(_02395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08301__S (.DIODE(_02395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08246__S0 (.DIODE(_02395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08208__S (.DIODE(_02395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08103__S (.DIODE(_02395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08046__S0 (.DIODE(_02395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07979__S0 (.DIODE(_02395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07957__S (.DIODE(_02395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08464__B1 (.DIODE(_02399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08419__B1 (.DIODE(_02399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08397__B1 (.DIODE(_02399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08304__B1 (.DIODE(_02399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08280__B1 (.DIODE(_02399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08211__B1 (.DIODE(_02399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08107__B1 (.DIODE(_02399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08082__B1 (.DIODE(_02399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08034__A (.DIODE(_02399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07961__B1 (.DIODE(_02399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08608__S1 (.DIODE(_02402_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08583__A (.DIODE(_02402_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08513__A (.DIODE(_02402_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08469__S1 (.DIODE(_02402_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08355__A (.DIODE(_02402_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08309__S1 (.DIODE(_02402_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08238__A (.DIODE(_02402_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08113__S1 (.DIODE(_02402_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08038__A (.DIODE(_02402_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07967__A (.DIODE(_02402_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08584__S (.DIODE(_02403_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08582__S (.DIODE(_02403_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08514__S (.DIODE(_02403_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08512__S (.DIODE(_02403_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08356__S (.DIODE(_02403_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08354__S (.DIODE(_02403_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08239__S (.DIODE(_02403_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08237__S (.DIODE(_02403_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08037__S (.DIODE(_02403_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07966__S (.DIODE(_02403_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08713__S0 (.DIODE(_02406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08712__S0 (.DIODE(_02406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08587__A1 (.DIODE(_02406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08517__A1 (.DIODE(_02406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08359__A1 (.DIODE(_02406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08242__A1 (.DIODE(_02406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08155__A (.DIODE(_02406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08039__S (.DIODE(_02406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08018__A (.DIODE(_02406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07969__S (.DIODE(_02406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08686__B1 (.DIODE(_02408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08664__B1 (.DIODE(_02408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08585__B1 (.DIODE(_02408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08515__B1 (.DIODE(_02408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08357__B1 (.DIODE(_02408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08240__B1 (.DIODE(_02408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08040__B1 (.DIODE(_02408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08015__A (.DIODE(_02408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07984__A (.DIODE(_02408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07971__B1 (.DIODE(_02408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08585__A1 (.DIODE(_02413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08515__A1 (.DIODE(_02413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08361__B2 (.DIODE(_02413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08357__A1 (.DIODE(_02413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08244__B2 (.DIODE(_02413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08240__A1 (.DIODE(_02413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08044__B2 (.DIODE(_02413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08040__A1 (.DIODE(_02413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08029__A (.DIODE(_02413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07977__B2 (.DIODE(_02413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08601__S (.DIODE(_02414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08531__S (.DIODE(_02414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08373__S (.DIODE(_02414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08256__S (.DIODE(_02414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08244__C1 (.DIODE(_02414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08117__A (.DIODE(_02414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08056__S (.DIODE(_02414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08044__C1 (.DIODE(_02414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07994__S (.DIODE(_02414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07977__C1 (.DIODE(_02414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08619__B1 (.DIODE(_02418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08593__A (.DIODE(_02418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08523__A (.DIODE(_02418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08480__B1 (.DIODE(_02418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08365__A (.DIODE(_02418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08320__B1 (.DIODE(_02418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08248__A (.DIODE(_02418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08127__B1 (.DIODE(_02418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08048__A (.DIODE(_02418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07982__A (.DIODE(_02418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08598__A1 (.DIODE(_02422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08564__B1 (.DIODE(_02422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08528__A1 (.DIODE(_02422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08504__B1 (.DIODE(_02422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08428__B1 (.DIODE(_02422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08370__A1 (.DIODE(_02422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08253__A1 (.DIODE(_02422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08112__A (.DIODE(_02422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08053__A1 (.DIODE(_02422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07989__A1 (.DIODE(_02422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08689__B1 (.DIODE(_02423_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08667__B1 (.DIODE(_02423_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08645__B1 (.DIODE(_02423_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08595__S1 (.DIODE(_02423_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08552__B1 (.DIODE(_02423_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08525__S1 (.DIODE(_02423_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08367__S1 (.DIODE(_02423_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08250__S1 (.DIODE(_02423_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08050__S1 (.DIODE(_02423_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07986__S1 (.DIODE(_02423_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08596__S0 (.DIODE(_02428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08529__S0 (.DIODE(_02428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08526__S0 (.DIODE(_02428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08371__S0 (.DIODE(_02428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08368__S0 (.DIODE(_02428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08254__S0 (.DIODE(_02428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08251__S0 (.DIODE(_02428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08054__S0 (.DIODE(_02428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08051__S0 (.DIODE(_02428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07992__S0 (.DIODE(_02428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08599__S1 (.DIODE(_02429_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08596__S1 (.DIODE(_02429_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08529__S1 (.DIODE(_02429_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08526__S1 (.DIODE(_02429_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08371__S1 (.DIODE(_02429_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08368__S1 (.DIODE(_02429_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08254__S1 (.DIODE(_02429_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08054__S1 (.DIODE(_02429_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07993__S1 (.DIODE(_02429_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07992__S1 (.DIODE(_02429_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08715__C1 (.DIODE(_02433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08627__A1 (.DIODE(_02433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08578__C1 (.DIODE(_02433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08488__A1 (.DIODE(_02433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08442__C1 (.DIODE(_02433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08328__A1 (.DIODE(_02433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08257__B1 (.DIODE(_02433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08135__A1 (.DIODE(_02433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08057__B1 (.DIODE(_02433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07996__B1 (.DIODE(_02433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07998__A1 (.DIODE(_02435_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08003__A2 (.DIODE(_02439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08621__B_N (.DIODE(_02445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08611__S0 (.DIODE(_02445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08482__B_N (.DIODE(_02445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08472__S0 (.DIODE(_02445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08322__B_N (.DIODE(_02445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08312__S0 (.DIODE(_02445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08143__A (.DIODE(_02445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08129__B_N (.DIODE(_02445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08116__S0 (.DIODE(_02445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08009__A (.DIODE(_02445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08676__S0 (.DIODE(_02446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08654__S0 (.DIODE(_02446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08632__S0 (.DIODE(_02446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08539__S0 (.DIODE(_02446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08498__S0 (.DIODE(_02446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08339__S0 (.DIODE(_02446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08223__S0 (.DIODE(_02446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08176__S0 (.DIODE(_02446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08151__S0 (.DIODE(_02446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08011__S0 (.DIODE(_02446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08676__S1 (.DIODE(_02447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08654__S1 (.DIODE(_02447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08632__S1 (.DIODE(_02447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08539__S1 (.DIODE(_02447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08339__S1 (.DIODE(_02447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08223__S1 (.DIODE(_02447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08176__S1 (.DIODE(_02447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08171__S1 (.DIODE(_02447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08151__S1 (.DIODE(_02447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08011__S1 (.DIODE(_02447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08681__S0 (.DIODE(_02449_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08659__S0 (.DIODE(_02449_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08637__S0 (.DIODE(_02449_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08544__S0 (.DIODE(_02449_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08499__S0 (.DIODE(_02449_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08340__S0 (.DIODE(_02449_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08224__S0 (.DIODE(_02449_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08177__S0 (.DIODE(_02449_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08152__S0 (.DIODE(_02449_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08014__S0 (.DIODE(_02449_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08681__S1 (.DIODE(_02450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08659__S1 (.DIODE(_02450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08637__S1 (.DIODE(_02450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08544__S1 (.DIODE(_02450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08498__S1 (.DIODE(_02450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08340__S1 (.DIODE(_02450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08224__S1 (.DIODE(_02450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08177__S1 (.DIODE(_02450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08152__S1 (.DIODE(_02450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08014__S1 (.DIODE(_02450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08631__S (.DIODE(_02452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08572__A (.DIODE(_02452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08500__S (.DIODE(_02452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08345__B1 (.DIODE(_02452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08341__S (.DIODE(_02452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08229__B1 (.DIODE(_02452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08225__S (.DIODE(_02452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08142__S (.DIODE(_02452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08024__B1 (.DIODE(_02452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08016__S (.DIODE(_02452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08687__A1 (.DIODE(_02454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08665__A1 (.DIODE(_02454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08643__A1 (.DIODE(_02454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08550__A1 (.DIODE(_02454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08502__A (.DIODE(_02454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08343__A (.DIODE(_02454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08227__A (.DIODE(_02454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08182__A1 (.DIODE(_02454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08159__A1 (.DIODE(_02454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08020__A (.DIODE(_02454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08563__S (.DIODE(_02455_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08561__S (.DIODE(_02455_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08501__S (.DIODE(_02455_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08427__S (.DIODE(_02455_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08425__S (.DIODE(_02455_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08342__S (.DIODE(_02455_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08232__S (.DIODE(_02455_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08226__S (.DIODE(_02455_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08028__S (.DIODE(_02455_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08019__S (.DIODE(_02455_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08708__S0 (.DIODE(_02458_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08704__S (.DIODE(_02458_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08685__S (.DIODE(_02458_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08663__S (.DIODE(_02458_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08641__S (.DIODE(_02458_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08623__S (.DIODE(_02458_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08484__S (.DIODE(_02458_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08324__S (.DIODE(_02458_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08131__S (.DIODE(_02458_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08022__A (.DIODE(_02458_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08458__S (.DIODE(_02459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08413__S (.DIODE(_02459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08395__S (.DIODE(_02459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08344__S (.DIODE(_02459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08298__S (.DIODE(_02459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08278__S (.DIODE(_02459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08228__S (.DIODE(_02459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08205__S (.DIODE(_02459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08079__S (.DIODE(_02459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08023__S (.DIODE(_02459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08629__S0 (.DIODE(_02462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08571__S0 (.DIODE(_02462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08536__S0 (.DIODE(_02462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08435__S0 (.DIODE(_02462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08231__A1 (.DIODE(_02462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08230__B_N (.DIODE(_02462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08168__S0 (.DIODE(_02462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08138__S0 (.DIODE(_02462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08027__A1 (.DIODE(_02462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08026__B_N (.DIODE(_02462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08564__A1 (.DIODE(_02466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08508__B2 (.DIODE(_02466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08432__B2 (.DIODE(_02466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08428__A1 (.DIODE(_02466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08396__B2 (.DIODE(_02466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08350__B2 (.DIODE(_02466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08279__B2 (.DIODE(_02466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08233__B2 (.DIODE(_02466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08081__B2 (.DIODE(_02466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08030__B2 (.DIODE(_02466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08609__B1 (.DIODE(_02468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08598__C1 (.DIODE(_02468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08528__C1 (.DIODE(_02468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08470__B1 (.DIODE(_02468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08370__C1 (.DIODE(_02468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08310__B1 (.DIODE(_02468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08253__C1 (.DIODE(_02468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08114__B1 (.DIODE(_02468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08053__C1 (.DIODE(_02468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08032__A (.DIODE(_02468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08679__B1 (.DIODE(_02469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08657__B1 (.DIODE(_02469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08635__B1 (.DIODE(_02469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08542__B1 (.DIODE(_02469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08509__B1 (.DIODE(_02469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08351__B1 (.DIODE(_02469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08234__C1 (.DIODE(_02469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08174__B1 (.DIODE(_02469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08148__B1 (.DIODE(_02469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08033__C1 (.DIODE(_02469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08693__C1 (.DIODE(_02471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08671__C1 (.DIODE(_02471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08649__C1 (.DIODE(_02471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08556__C1 (.DIODE(_02471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08510__C1 (.DIODE(_02471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08352__C1 (.DIODE(_02471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08235__C1 (.DIODE(_02471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08188__C1 (.DIODE(_02471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08166__C1 (.DIODE(_02471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08035__C1 (.DIODE(_02471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08036__C1 (.DIODE(_02472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08059__A1 (.DIODE(_02494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08691__B2 (.DIODE(_02508_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08669__B2 (.DIODE(_02508_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08647__B2 (.DIODE(_02508_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08568__B2 (.DIODE(_02508_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08554__B2 (.DIODE(_02508_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08391__A1 (.DIODE(_02508_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08274__A1 (.DIODE(_02508_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08186__B2 (.DIODE(_02508_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08164__B2 (.DIODE(_02508_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08075__A1 (.DIODE(_02508_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08470__A1 (.DIODE(_02515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08459__C1 (.DIODE(_02515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08414__C1 (.DIODE(_02515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08396__C1 (.DIODE(_02515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08310__A1 (.DIODE(_02515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08299__C1 (.DIODE(_02515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08279__C1 (.DIODE(_02515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08206__C1 (.DIODE(_02515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08114__A1 (.DIODE(_02515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08081__C1 (.DIODE(_02515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08083__B1 (.DIODE(_02517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08084__C1 (.DIODE(_02518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08494__S0 (.DIODE(_02523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08449__S0 (.DIODE(_02523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08404__S0 (.DIODE(_02523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08382__S0 (.DIODE(_02523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08335__S0 (.DIODE(_02523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08288__S0 (.DIODE(_02523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08265__S0 (.DIODE(_02523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08219__S0 (.DIODE(_02523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08196__S0 (.DIODE(_02523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08090__S0 (.DIODE(_02523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08496__S (.DIODE(_02526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08451__S (.DIODE(_02526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08406__S (.DIODE(_02526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08384__S (.DIODE(_02526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08337__S (.DIODE(_02526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08291__S (.DIODE(_02526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08267__S (.DIODE(_02526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08221__S (.DIODE(_02526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08198__S (.DIODE(_02526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08093__S (.DIODE(_02526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08701__C1 (.DIODE(_02538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08642__B1 (.DIODE(_02538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08549__B1 (.DIODE(_02538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08462__B1 (.DIODE(_02538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08417__B1 (.DIODE(_02538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08302__B1 (.DIODE(_02538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08209__B1 (.DIODE(_02538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08181__B1 (.DIODE(_02538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08158__B1 (.DIODE(_02538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08105__B1 (.DIODE(_02538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08109__C1 (.DIODE(_02542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09606__A2 (.DIODE(_02543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09425__A2 (.DIODE(_02543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09267__A2 (.DIODE(_02543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08945__A2 (.DIODE(_02543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08716__A (.DIODE(_02543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08628__A2 (.DIODE(_02543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08489__A2 (.DIODE(_02543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08443__B (.DIODE(_02543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08329__A2 (.DIODE(_02543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08136__A2 (.DIODE(_02543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08691__C1 (.DIODE(_02550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08669__C1 (.DIODE(_02550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08647__C1 (.DIODE(_02550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08568__C1 (.DIODE(_02550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08554__C1 (.DIODE(_02550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08473__S (.DIODE(_02550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08313__S (.DIODE(_02550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08186__C1 (.DIODE(_02550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08164__C1 (.DIODE(_02550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08118__S (.DIODE(_02550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08690__S (.DIODE(_02553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08668__S (.DIODE(_02553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08646__S (.DIODE(_02553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08567__S (.DIODE(_02553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08553__S (.DIODE(_02553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08431__S (.DIODE(_02553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08315__S0 (.DIODE(_02553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08185__S (.DIODE(_02553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08163__S (.DIODE(_02553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08121__S0 (.DIODE(_02553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08615__S1 (.DIODE(_02555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08614__S1 (.DIODE(_02555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08566__B1 (.DIODE(_02555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08476__S1 (.DIODE(_02555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08475__S1 (.DIODE(_02555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08430__B1 (.DIODE(_02555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08316__S1 (.DIODE(_02555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08184__B1 (.DIODE(_02555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08162__B1 (.DIODE(_02555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08123__S1 (.DIODE(_02555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08136__B1 (.DIODE(_02568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08680__A1 (.DIODE(_02569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08658__A1 (.DIODE(_02569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08636__A1 (.DIODE(_02569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08543__A1 (.DIODE(_02569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08497__B2 (.DIODE(_02569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08452__B2 (.DIODE(_02569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08407__B2 (.DIODE(_02569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08385__B2 (.DIODE(_02569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08175__A1 (.DIODE(_02569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08149__A1 (.DIODE(_02569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08674__S0 (.DIODE(_02571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08673__S0 (.DIODE(_02571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08652__S0 (.DIODE(_02571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08651__S0 (.DIODE(_02571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08630__S0 (.DIODE(_02571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08575__S0 (.DIODE(_02571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08537__S0 (.DIODE(_02571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08439__S0 (.DIODE(_02571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08169__S0 (.DIODE(_02571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08141__S0 (.DIODE(_02571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08674__S1 (.DIODE(_02572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08673__S1 (.DIODE(_02572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08652__S1 (.DIODE(_02572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08651__S1 (.DIODE(_02572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08630__S1 (.DIODE(_02572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08629__S1 (.DIODE(_02572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08537__S1 (.DIODE(_02572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08439__S1 (.DIODE(_02572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08169__S1 (.DIODE(_02572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08141__S1 (.DIODE(_02572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08492__S0 (.DIODE(_02575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08447__S0 (.DIODE(_02575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08402__S0 (.DIODE(_02575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08380__S0 (.DIODE(_02575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08333__S0 (.DIODE(_02575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08286__S0 (.DIODE(_02575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08263__S0 (.DIODE(_02575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08217__S0 (.DIODE(_02575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08171__S0 (.DIODE(_02575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08145__S0 (.DIODE(_02575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08492__S1 (.DIODE(_02576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08447__S1 (.DIODE(_02576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08402__S1 (.DIODE(_02576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08380__S1 (.DIODE(_02576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08333__S1 (.DIODE(_02576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08286__S1 (.DIODE(_02576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08263__S1 (.DIODE(_02576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08217__S1 (.DIODE(_02576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08194__S1 (.DIODE(_02576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08145__S1 (.DIODE(_02576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08693__A1 (.DIODE(_02582_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08671__A1 (.DIODE(_02582_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08649__A1 (.DIODE(_02582_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08556__A1 (.DIODE(_02582_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08510__A1 (.DIODE(_02582_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08434__A1 (.DIODE(_02582_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08352__A1 (.DIODE(_02582_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08235__A1 (.DIODE(_02582_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08188__A1 (.DIODE(_02582_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08166__A1 (.DIODE(_02582_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08670__A (.DIODE(_02586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08648__A (.DIODE(_02586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08555__A (.DIODE(_02586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08493__B1 (.DIODE(_02586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08448__B1 (.DIODE(_02586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08403__B1 (.DIODE(_02586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08381__B1 (.DIODE(_02586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08334__B1 (.DIODE(_02586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08187__A (.DIODE(_02586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08165__A (.DIODE(_02586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11164__A1 (.DIODE(_02587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08684__S (.DIODE(_02587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08662__S (.DIODE(_02587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08640__S (.DIODE(_02587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08547__S (.DIODE(_02587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08507__S (.DIODE(_02587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08503__S (.DIODE(_02587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08349__S (.DIODE(_02587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08179__S (.DIODE(_02587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08156__S (.DIODE(_02587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08644__B_N (.DIODE(_02592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08576__S0 (.DIODE(_02592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08566__A1 (.DIODE(_02592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08565__B_N (.DIODE(_02592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08551__B_N (.DIODE(_02592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08440__S0 (.DIODE(_02592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08430__A1 (.DIODE(_02592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08429__B_N (.DIODE(_02592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08183__B_N (.DIODE(_02592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08161__B_N (.DIODE(_02592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08189__B2 (.DIODE(_02606_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08189__C1 (.DIODE(_02619_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08491__A (.DIODE(_02620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08446__A (.DIODE(_02620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08436__A (.DIODE(_02620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08401__A (.DIODE(_02620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08379__A (.DIODE(_02620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08332__A (.DIODE(_02620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08285__A (.DIODE(_02620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08262__A (.DIODE(_02620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08216__A (.DIODE(_02620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08192__A (.DIODE(_02620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08540__A (.DIODE(_02623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08493__A1 (.DIODE(_02623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08448__A1 (.DIODE(_02623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08403__A1 (.DIODE(_02623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08381__A1 (.DIODE(_02623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08334__A1 (.DIODE(_02623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08287__A1 (.DIODE(_02623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08264__A1 (.DIODE(_02623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08218__A1 (.DIODE(_02623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08195__A1 (.DIODE(_02623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08213__C1 (.DIODE(_02642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08573__S1 (.DIODE(_02643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08490__S1 (.DIODE(_02643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08445__S1 (.DIODE(_02643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08437__S1 (.DIODE(_02643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08400__S1 (.DIODE(_02643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08378__S1 (.DIODE(_02643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08331__S1 (.DIODE(_02643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08284__S1 (.DIODE(_02643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08261__S1 (.DIODE(_02643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08215__S1 (.DIODE(_02643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08236__C1 (.DIODE(_02664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08259__A1 (.DIODE(_02686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08264__A2 (.DIODE(_02690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08282__B2 (.DIODE(_02695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08694__B1 (.DIODE(_02709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08672__B1 (.DIODE(_02709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08650__B1 (.DIODE(_02709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08557__B1 (.DIODE(_02709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08511__B1 (.DIODE(_02709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08466__B1 (.DIODE(_02709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08421__B1 (.DIODE(_02709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08399__B1 (.DIODE(_02709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08353__B1 (.DIODE(_02709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08306__B1 (.DIODE(_02709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08559__S1 (.DIODE(_02715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08558__S1 (.DIODE(_02715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08495__S1 (.DIODE(_02715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08450__S1 (.DIODE(_02715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08423__S1 (.DIODE(_02715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08422__S1 (.DIODE(_02715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08405__S1 (.DIODE(_02715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08383__S1 (.DIODE(_02715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08336__S1 (.DIODE(_02715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08290__S1 (.DIODE(_02715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08306__B2 (.DIODE(_02718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08306__C1 (.DIODE(_02731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08328__A2 (.DIODE(_02739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08329__B1 (.DIODE(_02753_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08993__A2 (.DIODE(_02754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08694__A2 (.DIODE(_02754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08672__A2 (.DIODE(_02754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08650__A2 (.DIODE(_02754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08557__A2 (.DIODE(_02754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08511__A2 (.DIODE(_02754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08466__A2 (.DIODE(_02754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08421__A2 (.DIODE(_02754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08399__A2 (.DIODE(_02754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08353__A2 (.DIODE(_02754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08353__B2 (.DIODE(_02762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08559__S0 (.DIODE(_02770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08558__S0 (.DIODE(_02770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08506__A1 (.DIODE(_02770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08505__B_N (.DIODE(_02770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08460__S (.DIODE(_02770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08423__S0 (.DIODE(_02770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08422__S0 (.DIODE(_02770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08415__S (.DIODE(_02770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08348__A1 (.DIODE(_02770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08347__B_N (.DIODE(_02770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08353__C1 (.DIODE(_02776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08376__A1 (.DIODE(_02798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08399__B2 (.DIODE(_02807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08399__C1 (.DIODE(_02820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08421__B2 (.DIODE(_02828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08421__C1 (.DIODE(_02841_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08444__A2 (.DIODE(_02854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08444__A3 (.DIODE(_02862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08466__B2 (.DIODE(_02871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08466__C1 (.DIODE(_02884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08487__A2 (.DIODE(_02895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08489__B1 (.DIODE(_02906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08511__B2 (.DIODE(_02914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08511__C1 (.DIODE(_02927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08534__A1 (.DIODE(_02949_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08557__B2 (.DIODE(_02958_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08557__C1 (.DIODE(_02971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08581__A2 (.DIODE(_02984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08581__A3 (.DIODE(_02992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09719__A2 (.DIODE(_02993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09674__A2 (.DIODE(_02993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09628__A2 (.DIODE(_02993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09583__A2 (.DIODE(_02993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09561__A2 (.DIODE(_02993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09515__A2 (.DIODE(_02993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09379__B (.DIODE(_02993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09115__B (.DIODE(_02993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09038__B (.DIODE(_02993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08580__B (.DIODE(_02993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08604__A1 (.DIODE(_03016_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08628__B1 (.DIODE(_03039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08650__B2 (.DIODE(_03047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08650__C1 (.DIODE(_03060_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08672__B2 (.DIODE(_03068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08672__C1 (.DIODE(_03081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08694__B2 (.DIODE(_03089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08694__C1 (.DIODE(_03102_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08716__C_N (.DIODE(_03123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08717__B1 (.DIODE(_03124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09695__C1 (.DIODE(_03233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09605__A1 (.DIODE(_03233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09424__A1 (.DIODE(_03233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09378__C1 (.DIODE(_03233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09266__A1 (.DIODE(_03233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09114__C1 (.DIODE(_03233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09066__B1 (.DIODE(_03233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09037__C1 (.DIODE(_03233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08990__A (.DIODE(_03233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08944__A1 (.DIODE(_03233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09632__B1 (.DIODE(_03235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09519__B1 (.DIODE(_03235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09473__B1 (.DIODE(_03235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09293__B1 (.DIODE(_03235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09171__B1 (.DIODE(_03235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09120__B1 (.DIODE(_03235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09055__A (.DIODE(_03235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09053__A (.DIODE(_03235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09043__B1 (.DIODE(_03235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08894__A (.DIODE(_03235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09681__B1 (.DIODE(_03236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09645__A1 (.DIODE(_03236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09532__A1 (.DIODE(_03236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09486__A1 (.DIODE(_03236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09364__B1 (.DIODE(_03236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09306__A1 (.DIODE(_03236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09184__A1 (.DIODE(_03236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09100__B1 (.DIODE(_03236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09008__B1 (.DIODE(_03236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08900__A (.DIODE(_03236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09647__S0 (.DIODE(_03237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09534__S0 (.DIODE(_03237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09488__S0 (.DIODE(_03237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09308__S0 (.DIODE(_03237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09186__S0 (.DIODE(_03237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09135__S0 (.DIODE(_03237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09064__S0 (.DIODE(_03237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08935__A (.DIODE(_03237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08907__A (.DIODE(_03237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08896__A (.DIODE(_03237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09642__S0 (.DIODE(_03238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09586__S0 (.DIODE(_03238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09529__S0 (.DIODE(_03238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09483__S0 (.DIODE(_03238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09405__S0 (.DIODE(_03238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09247__S0 (.DIODE(_03238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09245__S0 (.DIODE(_03238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09201__A (.DIODE(_03238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08905__S0 (.DIODE(_03238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08899__S0 (.DIODE(_03238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10779__B2 (.DIODE(_03239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09647__S1 (.DIODE(_03239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09534__S1 (.DIODE(_03239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09488__S1 (.DIODE(_03239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09308__S1 (.DIODE(_03239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09295__B1 (.DIODE(_03239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09173__B1 (.DIODE(_03239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09122__B1 (.DIODE(_03239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09046__B1 (.DIODE(_03239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08898__A (.DIODE(_03239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09630__A (.DIODE(_03240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09584__S1 (.DIODE(_03240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09517__A (.DIODE(_03240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09403__S1 (.DIODE(_03240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09245__S1 (.DIODE(_03240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09223__A (.DIODE(_03240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09153__A (.DIODE(_03240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09150__A (.DIODE(_03240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08954__A (.DIODE(_03240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08899__S1 (.DIODE(_03240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09602__C1 (.DIODE(_03243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09590__S (.DIODE(_03243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09421__C1 (.DIODE(_03243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09409__S (.DIODE(_03243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09263__C1 (.DIODE(_03243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09034__A (.DIODE(_03243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08999__A (.DIODE(_03243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08966__A (.DIODE(_03243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08941__C1 (.DIODE(_03243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08902__A (.DIODE(_03243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09712__C1 (.DIODE(_03244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09587__A1 (.DIODE(_03244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09406__A1 (.DIODE(_03244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09354__C1 (.DIODE(_03244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09328__C1 (.DIODE(_03244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09282__C1 (.DIODE(_03244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09248__A1 (.DIODE(_03244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09090__C1 (.DIODE(_03244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08989__C1 (.DIODE(_03244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08906__A1 (.DIODE(_03244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09643__S1 (.DIODE(_03245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09530__S1 (.DIODE(_03245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09484__S1 (.DIODE(_03245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09304__S1 (.DIODE(_03245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09182__S1 (.DIODE(_03245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09131__S1 (.DIODE(_03245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09058__S1 (.DIODE(_03245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09056__A (.DIODE(_03245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09012__A (.DIODE(_03245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08904__A (.DIODE(_03245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09586__S1 (.DIODE(_03246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09471__A (.DIODE(_03246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09405__S1 (.DIODE(_03246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09291__A (.DIODE(_03246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09247__S1 (.DIODE(_03246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09169__A (.DIODE(_03246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09118__A (.DIODE(_03246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09080__A (.DIODE(_03246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09041__A (.DIODE(_03246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08905__S1 (.DIODE(_03246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09588__S0 (.DIODE(_03249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09584__S0 (.DIODE(_03249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09408__S0 (.DIODE(_03249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09407__S0 (.DIODE(_03249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09403__S0 (.DIODE(_03249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09250__S0 (.DIODE(_03249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09249__S0 (.DIODE(_03249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08953__A (.DIODE(_03249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08911__S0 (.DIODE(_03249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08910__S0 (.DIODE(_03249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09634__B1 (.DIODE(_03250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09521__B1 (.DIODE(_03250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09480__S1 (.DIODE(_03250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09475__B1 (.DIODE(_03250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09300__S1 (.DIODE(_03250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09178__S1 (.DIODE(_03250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09127__S1 (.DIODE(_03250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09052__S1 (.DIODE(_03250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08963__A (.DIODE(_03250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08909__A (.DIODE(_03250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09589__S1 (.DIODE(_03251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09588__S1 (.DIODE(_03251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09408__S1 (.DIODE(_03251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09407__S1 (.DIODE(_03251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09250__S1 (.DIODE(_03251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09249__S1 (.DIODE(_03251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08960__A (.DIODE(_03251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08950__A (.DIODE(_03251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08911__S1 (.DIODE(_03251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08910__S1 (.DIODE(_03251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09648__S (.DIODE(_03254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09535__S (.DIODE(_03254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09489__S (.DIODE(_03254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09309__S (.DIODE(_03254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09187__S (.DIODE(_03254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09175__C1 (.DIODE(_03254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09136__S (.DIODE(_03254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09124__C1 (.DIODE(_03254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09049__C1 (.DIODE(_03254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08913__A (.DIODE(_03254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09671__C1 (.DIODE(_03255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09625__C1 (.DIODE(_03255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09580__C1 (.DIODE(_03255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09558__C1 (.DIODE(_03255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09466__C1 (.DIODE(_03255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09444__C1 (.DIODE(_03255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09399__C1 (.DIODE(_03255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09251__S (.DIODE(_03255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09026__A (.DIODE(_03255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08914__S (.DIODE(_03255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09649__A1 (.DIODE(_03258_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09641__C1 (.DIODE(_03258_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09528__C1 (.DIODE(_03258_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09482__C1 (.DIODE(_03258_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09302__C1 (.DIODE(_03258_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09180__C1 (.DIODE(_03258_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09129__C1 (.DIODE(_03258_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09054__C1 (.DIODE(_03258_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08968__A (.DIODE(_03258_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08917__A (.DIODE(_03258_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09695__B2 (.DIODE(_03259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09604__A1 (.DIODE(_03259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09423__A1 (.DIODE(_03259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09410__B2 (.DIODE(_03259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09378__B2 (.DIODE(_03259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09265__A1 (.DIODE(_03259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09252__B2 (.DIODE(_03259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08971__A (.DIODE(_03259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08943__A1 (.DIODE(_03259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08918__B2 (.DIODE(_03259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09670__S (.DIODE(_03261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09624__S (.DIODE(_03261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09579__S (.DIODE(_03261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09557__S (.DIODE(_03261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09465__S (.DIODE(_03261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09443__S (.DIODE(_03261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09411__S0 (.DIODE(_03261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09398__S (.DIODE(_03261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09253__S0 (.DIODE(_03261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08921__S0 (.DIODE(_03261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09592__S1 (.DIODE(_03262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09510__B1 (.DIODE(_03262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09412__S1 (.DIODE(_03262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09411__S1 (.DIODE(_03262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09254__S1 (.DIODE(_03262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09253__S1 (.DIODE(_03262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09161__B1 (.DIODE(_03262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08972__A (.DIODE(_03262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08922__S1 (.DIODE(_03262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08921__S1 (.DIODE(_03262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09637__C1 (.DIODE(_03266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09524__C1 (.DIODE(_03266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09478__C1 (.DIODE(_03266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09298__C1 (.DIODE(_03266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09176__C1 (.DIODE(_03266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09125__C1 (.DIODE(_03266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09050__C1 (.DIODE(_03266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09028__A (.DIODE(_03266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08956__A (.DIODE(_03266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08925__A (.DIODE(_03266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09691__B1 (.DIODE(_03267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09603__A1 (.DIODE(_03267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09422__A1 (.DIODE(_03267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09374__B1 (.DIODE(_03267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09264__A1 (.DIODE(_03267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09184__C1 (.DIODE(_03267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09133__C1 (.DIODE(_03267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09110__B1 (.DIODE(_03267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09060__C1 (.DIODE(_03267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08942__A1 (.DIODE(_03267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09688__S1 (.DIODE(_03268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09598__A1 (.DIODE(_03268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09417__A1 (.DIODE(_03268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09381__S1 (.DIODE(_03268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09371__S1 (.DIODE(_03268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09259__A1 (.DIODE(_03268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09217__S1 (.DIODE(_03268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09107__S1 (.DIODE(_03268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09024__S1 (.DIODE(_03268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08934__A1 (.DIODE(_03268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09596__S (.DIODE(_03269_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09415__S (.DIODE(_03269_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09300__S0 (.DIODE(_03269_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09257__S (.DIODE(_03269_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09178__S0 (.DIODE(_03269_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09127__S0 (.DIODE(_03269_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09052__S0 (.DIODE(_03269_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08948__A (.DIODE(_03269_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08931__S (.DIODE(_03269_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08928__A (.DIODE(_03269_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09714__S (.DIODE(_03270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09638__S0 (.DIODE(_03270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09525__S0 (.DIODE(_03270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09479__S0 (.DIODE(_03270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09299__S0 (.DIODE(_03270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09256__S (.DIODE(_03270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09177__S0 (.DIODE(_03270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09126__S0 (.DIODE(_03270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09051__S0 (.DIODE(_03270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08929__S (.DIODE(_03270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09636__B2 (.DIODE(_03272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09597__A1 (.DIODE(_03272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09523__B2 (.DIODE(_03272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09416__A1 (.DIODE(_03272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09258__A1 (.DIODE(_03272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09210__A (.DIODE(_03272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09015__A (.DIODE(_03272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08979__A (.DIODE(_03272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08940__A (.DIODE(_03272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08933__A1 (.DIODE(_03272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09640__A (.DIODE(_03274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09597__B1 (.DIODE(_03274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09527__A (.DIODE(_03274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09481__A (.DIODE(_03274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09416__B1 (.DIODE(_03274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09301__A (.DIODE(_03274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09258__B1 (.DIODE(_03274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09179__A (.DIODE(_03274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09128__A (.DIODE(_03274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08933__B1 (.DIODE(_03274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09599__B_N (.DIODE(_03277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09589__S0 (.DIODE(_03277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09418__B_N (.DIODE(_03277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09260__B_N (.DIODE(_03277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09222__A (.DIODE(_03277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09152__A (.DIODE(_03277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09149__A (.DIODE(_03277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08983__A (.DIODE(_03277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08937__A1 (.DIODE(_03277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08936__B_N (.DIODE(_03277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09665__S (.DIODE(_03280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09601__S (.DIODE(_03280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09420__S (.DIODE(_03280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09294__B_N (.DIODE(_03280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09262__S (.DIODE(_03280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09172__B_N (.DIODE(_03280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09121__B_N (.DIODE(_03280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09044__B_N (.DIODE(_03280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08986__A (.DIODE(_03280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08939__S (.DIODE(_03280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09666__A1 (.DIODE(_03282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09620__A1 (.DIODE(_03282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09602__B2 (.DIODE(_03282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09421__B2 (.DIODE(_03282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09263__B2 (.DIODE(_03282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09171__A1 (.DIODE(_03282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09120__A1 (.DIODE(_03282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09043__A1 (.DIODE(_03282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08988__A (.DIODE(_03282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08941__B2 (.DIODE(_03282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08945__B1 (.DIODE(_03286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09585__A (.DIODE(_03287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09404__A (.DIODE(_03287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09349__B1 (.DIODE(_03287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09285__B1 (.DIODE(_03287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09246__A (.DIODE(_03287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09212__B1 (.DIODE(_03287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09085__B1 (.DIODE(_03287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09022__A (.DIODE(_03287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08981__B1 (.DIODE(_03287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08947__A (.DIODE(_03287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09708__S (.DIODE(_03288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09657__A (.DIODE(_03288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09611__A (.DIODE(_03288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09566__A (.DIODE(_03288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09544__A (.DIODE(_03288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09452__A (.DIODE(_03288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09430__A (.DIODE(_03288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09385__A (.DIODE(_03288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09225__A (.DIODE(_03288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08952__A (.DIODE(_03288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09600__A1 (.DIODE(_03289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09419__A1 (.DIODE(_03289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09348__S (.DIODE(_03289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09330__S (.DIODE(_03289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09284__S (.DIODE(_03289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09261__A1 (.DIODE(_03289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09211__S (.DIODE(_03289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09084__S (.DIODE(_03289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08980__S (.DIODE(_03289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08949__A (.DIODE(_03289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09352__A1 (.DIODE(_03290_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09351__B_N (.DIODE(_03290_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09314__S0 (.DIODE(_03290_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09268__S0 (.DIODE(_03290_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09192__S0 (.DIODE(_03290_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09141__S0 (.DIODE(_03290_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09088__A1 (.DIODE(_03290_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09071__S0 (.DIODE(_03290_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08985__A1 (.DIODE(_03290_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08951__S0 (.DIODE(_03290_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09698__S1 (.DIODE(_03291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09662__S1 (.DIODE(_03291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09494__S1 (.DIODE(_03291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09336__S1 (.DIODE(_03291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09314__S1 (.DIODE(_03291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09268__S1 (.DIODE(_03291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09192__S1 (.DIODE(_03291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09141__S1 (.DIODE(_03291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09071__S1 (.DIODE(_03291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08951__S1 (.DIODE(_03291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09658__S0 (.DIODE(_03294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09612__S0 (.DIODE(_03294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09567__S0 (.DIODE(_03294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09338__S0 (.DIODE(_03294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09316__S0 (.DIODE(_03294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09270__S0 (.DIODE(_03294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09194__S0 (.DIODE(_03294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09143__S0 (.DIODE(_03294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09073__S0 (.DIODE(_03294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08955__S0 (.DIODE(_03294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09658__S1 (.DIODE(_03295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09612__S1 (.DIODE(_03295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09567__S1 (.DIODE(_03295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09545__S1 (.DIODE(_03295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09316__S1 (.DIODE(_03295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09270__S1 (.DIODE(_03295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09194__S1 (.DIODE(_03295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09143__S1 (.DIODE(_03295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09073__S1 (.DIODE(_03295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08955__S1 (.DIODE(_03295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09686__C1 (.DIODE(_03297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09497__B1 (.DIODE(_03297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09369__C1 (.DIODE(_03297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09339__B1 (.DIODE(_03297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09317__B1 (.DIODE(_03297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09271__B1 (.DIODE(_03297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09195__B1 (.DIODE(_03297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09144__B1 (.DIODE(_03297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09074__B1 (.DIODE(_03297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08957__B1 (.DIODE(_03297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10770__B2 (.DIODE(_03299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09595__S (.DIODE(_03299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09414__S (.DIODE(_03299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09218__A (.DIODE(_03299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09030__A (.DIODE(_03299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09023__A (.DIODE(_03299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08995__A (.DIODE(_03299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08977__A (.DIODE(_03299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08962__A (.DIODE(_03299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08959__A (.DIODE(_03299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09698__S0 (.DIODE(_03300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09690__S0 (.DIODE(_03300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09494__S0 (.DIODE(_03300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09373__S0 (.DIODE(_03300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09336__S0 (.DIODE(_03300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09145__S0 (.DIODE(_03300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09109__S0 (.DIODE(_03300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09075__S0 (.DIODE(_03300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09027__S0 (.DIODE(_03300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08961__S0 (.DIODE(_03300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09690__S1 (.DIODE(_03301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09373__S1 (.DIODE(_03301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09318__S1 (.DIODE(_03301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09272__S1 (.DIODE(_03301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09196__S1 (.DIODE(_03301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09145__S1 (.DIODE(_03301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09109__S1 (.DIODE(_03301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09075__S1 (.DIODE(_03301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09027__S1 (.DIODE(_03301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08961__S1 (.DIODE(_03301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09702__S0 (.DIODE(_03303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09498__S0 (.DIODE(_03303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09340__S0 (.DIODE(_03303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09318__S0 (.DIODE(_03303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09272__S0 (.DIODE(_03303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09197__S0 (.DIODE(_03303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09196__S0 (.DIODE(_03303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09146__S0 (.DIODE(_03303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09076__S0 (.DIODE(_03303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08965__S0 (.DIODE(_03303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09638__S1 (.DIODE(_03304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09525__S1 (.DIODE(_03304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09479__S1 (.DIODE(_03304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09299__S1 (.DIODE(_03304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09177__S1 (.DIODE(_03304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09126__S1 (.DIODE(_03304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09051__S1 (.DIODE(_03304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09001__A (.DIODE(_03304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08996__A (.DIODE(_03304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08964__A (.DIODE(_03304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09702__S1 (.DIODE(_03305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09498__S1 (.DIODE(_03305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09341__S1 (.DIODE(_03305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09340__S1 (.DIODE(_03305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09319__S1 (.DIODE(_03305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09273__S1 (.DIODE(_03305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09197__S1 (.DIODE(_03305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09146__S1 (.DIODE(_03305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09076__S1 (.DIODE(_03305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08965__S1 (.DIODE(_03305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09663__S (.DIODE(_03307_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09617__S (.DIODE(_03307_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09572__S (.DIODE(_03307_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09550__S (.DIODE(_03307_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09458__S (.DIODE(_03307_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09436__S (.DIODE(_03307_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09198__S (.DIODE(_03307_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09147__S (.DIODE(_03307_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09077__S (.DIODE(_03307_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08967__S (.DIODE(_03307_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09591__B2 (.DIODE(_03309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09536__A1 (.DIODE(_03309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09490__A1 (.DIODE(_03309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09310__A1 (.DIODE(_03309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09188__A1 (.DIODE(_03309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09137__A1 (.DIODE(_03309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09066__A1 (.DIODE(_03309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09036__A (.DIODE(_03309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08994__A (.DIODE(_03309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08969__A (.DIODE(_03309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09705__B2 (.DIODE(_03310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09687__A1 (.DIODE(_03310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09501__B2 (.DIODE(_03310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09343__B2 (.DIODE(_03310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09321__B2 (.DIODE(_03310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09275__B2 (.DIODE(_03310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09199__B2 (.DIODE(_03310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09148__B2 (.DIODE(_03310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09078__B2 (.DIODE(_03310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08970__B2 (.DIODE(_03310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08993__B2 (.DIODE(_03311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09718__A1 (.DIODE(_03312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09401__A1 (.DIODE(_03312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09356__A1 (.DIODE(_03312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09334__A1 (.DIODE(_03312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09288__A1 (.DIODE(_03312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09243__A1 (.DIODE(_03312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09215__A1 (.DIODE(_03312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09166__A1 (.DIODE(_03312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09092__A1 (.DIODE(_03312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08992__A1 (.DIODE(_03312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09706__S1 (.DIODE(_03313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09679__A (.DIODE(_03313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09362__A (.DIODE(_03313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09344__S1 (.DIODE(_03313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09322__S1 (.DIODE(_03313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09276__S1 (.DIODE(_03313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09200__S1 (.DIODE(_03313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09079__S1 (.DIODE(_03313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08974__S1 (.DIODE(_03313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08973__S1 (.DIODE(_03313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09701__A1 (.DIODE(_03316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09497__A1 (.DIODE(_03316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09339__A1 (.DIODE(_03316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09317__A1 (.DIODE(_03316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09271__A1 (.DIODE(_03316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09195__A1 (.DIODE(_03316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09144__A1 (.DIODE(_03316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09082__S (.DIODE(_03316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09074__A1 (.DIODE(_03316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08976__S (.DIODE(_03316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09703__S0 (.DIODE(_03318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09499__S0 (.DIODE(_03318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09347__S (.DIODE(_03318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09341__S0 (.DIODE(_03318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09319__S0 (.DIODE(_03318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09283__S (.DIODE(_03318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09273__S0 (.DIODE(_03318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09209__S (.DIODE(_03318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09083__S (.DIODE(_03318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08978__S (.DIODE(_03318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09671__B2 (.DIODE(_03320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09625__B2 (.DIODE(_03320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09580__B2 (.DIODE(_03320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09558__B2 (.DIODE(_03320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09466__B2 (.DIODE(_03320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09444__B2 (.DIODE(_03320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09399__B2 (.DIODE(_03320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09349__A1 (.DIODE(_03320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09085__A1 (.DIODE(_03320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08981__A1 (.DIODE(_03320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09710__A1 (.DIODE(_03324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09709__B_N (.DIODE(_03324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09326__A1 (.DIODE(_03324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09325__B_N (.DIODE(_03324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09280__A1 (.DIODE(_03324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09279__B_N (.DIODE(_03324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09205__A1 (.DIODE(_03324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09204__B_N (.DIODE(_03324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09087__B_N (.DIODE(_03324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08984__B_N (.DIODE(_03324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09551__S (.DIODE(_03327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09507__S (.DIODE(_03327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09459__S (.DIODE(_03327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09437__S (.DIODE(_03327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09392__S (.DIODE(_03327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09353__S (.DIODE(_03327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09232__S (.DIODE(_03327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09158__S (.DIODE(_03327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09089__S (.DIODE(_03327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08987__S (.DIODE(_03327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09712__B2 (.DIODE(_03329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09508__A1 (.DIODE(_03329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09354__B2 (.DIODE(_03329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09328__B2 (.DIODE(_03329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09282__B2 (.DIODE(_03329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09208__B2 (.DIODE(_03329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09159__A1 (.DIODE(_03329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09090__B2 (.DIODE(_03329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09008__A1 (.DIODE(_03329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08989__B2 (.DIODE(_03329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09717__B1 (.DIODE(_03331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09355__B1 (.DIODE(_03331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09333__B1 (.DIODE(_03331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09287__B1 (.DIODE(_03331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09214__B1 (.DIODE(_03331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09165__A (.DIODE(_03331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09091__B1 (.DIODE(_03331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08991__B1 (.DIODE(_03331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09673__A1 (.DIODE(_03334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09627__A1 (.DIODE(_03334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09582__A1 (.DIODE(_03334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09560__A1 (.DIODE(_03334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09514__A1 (.DIODE(_03334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09468__A1 (.DIODE(_03334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09446__A1 (.DIODE(_03334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09370__A1 (.DIODE(_03334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09106__A1 (.DIODE(_03334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09021__A1 (.DIODE(_03334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09713__S (.DIODE(_03335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09676__S0 (.DIODE(_03335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09675__S0 (.DIODE(_03335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09359__S0 (.DIODE(_03335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09358__S0 (.DIODE(_03335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09329__S (.DIODE(_03335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09095__S0 (.DIODE(_03335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09094__S0 (.DIODE(_03335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08998__S0 (.DIODE(_03335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08997__S0 (.DIODE(_03335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09703__S1 (.DIODE(_03336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09676__S1 (.DIODE(_03336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09675__S1 (.DIODE(_03336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09499__S1 (.DIODE(_03336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09359__S1 (.DIODE(_03336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09358__S1 (.DIODE(_03336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09095__S1 (.DIODE(_03336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09094__S1 (.DIODE(_03336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08998__S1 (.DIODE(_03336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08997__S1 (.DIODE(_03336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09704__S (.DIODE(_03339_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09677__S (.DIODE(_03339_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09500__S (.DIODE(_03339_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09360__S (.DIODE(_03339_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09342__S (.DIODE(_03339_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09320__S (.DIODE(_03339_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09274__S (.DIODE(_03339_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09221__S (.DIODE(_03339_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09096__S (.DIODE(_03339_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09000__S (.DIODE(_03339_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09667__A1 (.DIODE(_03341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09621__A1 (.DIODE(_03341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09576__A1 (.DIODE(_03341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09554__A1 (.DIODE(_03341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09506__A (.DIODE(_03341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09462__A1 (.DIODE(_03341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09440__A1 (.DIODE(_03341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09157__A (.DIODE(_03341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09098__A (.DIODE(_03341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09005__A (.DIODE(_03341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09631__S (.DIODE(_03342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09518__S (.DIODE(_03342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09472__S (.DIODE(_03342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09292__S (.DIODE(_03342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09170__S (.DIODE(_03342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09119__S (.DIODE(_03342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09042__S (.DIODE(_03342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09040__S (.DIODE(_03342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09006__A (.DIODE(_03342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09003__A (.DIODE(_03342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09684__S (.DIODE(_03343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09678__S (.DIODE(_03343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09511__S (.DIODE(_03343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09367__S (.DIODE(_03343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09361__S (.DIODE(_03343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09240__S (.DIODE(_03343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09103__S (.DIODE(_03343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09097__S (.DIODE(_03343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09014__S (.DIODE(_03343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09004__S (.DIODE(_03343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09680__S (.DIODE(_03346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09664__S (.DIODE(_03346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09618__S (.DIODE(_03346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09573__S (.DIODE(_03346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09505__S (.DIODE(_03346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09363__S (.DIODE(_03346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09162__S (.DIODE(_03346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09156__S (.DIODE(_03346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09099__S (.DIODE(_03346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09007__S (.DIODE(_03346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09619__S (.DIODE(_03349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09574__S (.DIODE(_03349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09552__S (.DIODE(_03349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09460__S (.DIODE(_03349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09438__S (.DIODE(_03349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09393__S (.DIODE(_03349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09237__A (.DIODE(_03349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09233__S (.DIODE(_03349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09206__A (.DIODE(_03349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09010__A (.DIODE(_03349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09693__S0 (.DIODE(_03350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09683__A1 (.DIODE(_03350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09682__B_N (.DIODE(_03350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09376__S0 (.DIODE(_03350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09366__A1 (.DIODE(_03350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09365__B_N (.DIODE(_03350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09102__A1 (.DIODE(_03350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09101__B_N (.DIODE(_03350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09013__A1 (.DIODE(_03350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09011__B_N (.DIODE(_03350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09683__B1 (.DIODE(_03352_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09593__S1 (.DIODE(_03352_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09556__B1 (.DIODE(_03352_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09464__B1 (.DIODE(_03352_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09442__B1 (.DIODE(_03352_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09397__B1 (.DIODE(_03352_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09366__B1 (.DIODE(_03352_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09239__B1 (.DIODE(_03352_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09102__B1 (.DIODE(_03352_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09013__B1 (.DIODE(_03352_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09632__A1 (.DIODE(_03355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09519__A1 (.DIODE(_03355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09477__B2 (.DIODE(_03355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09473__A1 (.DIODE(_03355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09297__B2 (.DIODE(_03355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09293__A1 (.DIODE(_03355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09175__B2 (.DIODE(_03355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09124__B2 (.DIODE(_03355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09049__B2 (.DIODE(_03355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09016__A (.DIODE(_03355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09685__B2 (.DIODE(_03356_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09681__A1 (.DIODE(_03356_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09512__B2 (.DIODE(_03356_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09368__B2 (.DIODE(_03356_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09364__A1 (.DIODE(_03356_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09241__B2 (.DIODE(_03356_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09163__B2 (.DIODE(_03356_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09104__B2 (.DIODE(_03356_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09100__A1 (.DIODE(_03356_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09018__B2 (.DIODE(_03356_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09685__C1 (.DIODE(_03357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09641__A1 (.DIODE(_03357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09528__A1 (.DIODE(_03357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09482__A1 (.DIODE(_03357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09368__C1 (.DIODE(_03357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09302__A1 (.DIODE(_03357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09241__C1 (.DIODE(_03357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09180__A1 (.DIODE(_03357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09104__C1 (.DIODE(_03357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09018__C1 (.DIODE(_03357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09659__B1 (.DIODE(_03359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09613__B1 (.DIODE(_03359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09568__B1 (.DIODE(_03359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09546__B1 (.DIODE(_03359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09454__B1 (.DIODE(_03359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09432__B1 (.DIODE(_03359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09387__B1 (.DIODE(_03359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09227__B1 (.DIODE(_03359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09105__C1 (.DIODE(_03359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09020__C1 (.DIODE(_03359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09039__A2 (.DIODE(_03361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09699__A (.DIODE(_03362_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09495__A (.DIODE(_03362_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09337__A (.DIODE(_03362_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09315__A (.DIODE(_03362_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09269__A (.DIODE(_03362_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09193__A (.DIODE(_03362_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09142__A (.DIODE(_03362_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09108__A (.DIODE(_03362_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09072__A (.DIODE(_03362_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09025__A (.DIODE(_03362_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09688__S0 (.DIODE(_03363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09510__A1 (.DIODE(_03363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09509__B_N (.DIODE(_03363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09381__S0 (.DIODE(_03363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09371__S0 (.DIODE(_03363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09217__S0 (.DIODE(_03363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09161__A1 (.DIODE(_03363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09160__B_N (.DIODE(_03363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09107__S0 (.DIODE(_03363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09024__S0 (.DIODE(_03363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09691__A1 (.DIODE(_03366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09391__S (.DIODE(_03366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09374__A1 (.DIODE(_03366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09346__S (.DIODE(_03366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09324__S (.DIODE(_03366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09278__S (.DIODE(_03366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09231__S (.DIODE(_03366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09203__S (.DIODE(_03366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09110__A1 (.DIODE(_03366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09029__A1 (.DIODE(_03366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09701__B1 (.DIODE(_03368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09672__A (.DIODE(_03368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09626__A (.DIODE(_03368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09581__A (.DIODE(_03368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09559__A (.DIODE(_03368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09467__A (.DIODE(_03368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09445__A (.DIODE(_03368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09400__A (.DIODE(_03368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09242__A (.DIODE(_03368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09029__B1 (.DIODE(_03368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09037__A2 (.DIODE(_03369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09692__S0 (.DIODE(_03370_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09654__S0 (.DIODE(_03370_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09608__S0 (.DIODE(_03370_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09563__S0 (.DIODE(_03370_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09541__S0 (.DIODE(_03370_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09375__S0 (.DIODE(_03370_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09112__S0 (.DIODE(_03370_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09111__S0 (.DIODE(_03370_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09033__S0 (.DIODE(_03370_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09032__S0 (.DIODE(_03370_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09692__S1 (.DIODE(_03371_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09654__S1 (.DIODE(_03371_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09608__S1 (.DIODE(_03371_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09563__S1 (.DIODE(_03371_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09541__S1 (.DIODE(_03371_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09375__S1 (.DIODE(_03371_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09112__S1 (.DIODE(_03371_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09111__S1 (.DIODE(_03371_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09033__S1 (.DIODE(_03371_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09032__S1 (.DIODE(_03371_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09694__S (.DIODE(_03374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09655__S (.DIODE(_03374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09564__S (.DIODE(_03374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09542__S (.DIODE(_03374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09428__S (.DIODE(_03374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09383__S (.DIODE(_03374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09377__S (.DIODE(_03374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09208__C1 (.DIODE(_03374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09113__S (.DIODE(_03374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09035__S (.DIODE(_03374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09660__A1 (.DIODE(_03376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09614__A1 (.DIODE(_03376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09569__A1 (.DIODE(_03376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09547__A1 (.DIODE(_03376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09455__A1 (.DIODE(_03376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09433__A1 (.DIODE(_03376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09388__A1 (.DIODE(_03376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09228__A1 (.DIODE(_03376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09114__B2 (.DIODE(_03376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09037__B2 (.DIODE(_03376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09634__A1 (.DIODE(_03384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09633__B_N (.DIODE(_03384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09521__A1 (.DIODE(_03384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09520__B_N (.DIODE(_03384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09475__A1 (.DIODE(_03384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09474__B_N (.DIODE(_03384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09295__A1 (.DIODE(_03384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09173__A1 (.DIODE(_03384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09122__A1 (.DIODE(_03384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09046__A1 (.DIODE(_03384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11348__A1 (.DIODE(_03386_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09629__S (.DIODE(_03386_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09516__S (.DIODE(_03386_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09470__S (.DIODE(_03386_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09290__S (.DIODE(_03386_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09174__S (.DIODE(_03386_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09168__S (.DIODE(_03386_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09123__S (.DIODE(_03386_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09117__S (.DIODE(_03386_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09048__S (.DIODE(_03386_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09689__A (.DIODE(_03394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09609__S (.DIODE(_03394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09508__B1 (.DIODE(_03394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09504__S (.DIODE(_03394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09450__S (.DIODE(_03394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09372__A (.DIODE(_03394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09159__B1 (.DIODE(_03394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09155__S (.DIODE(_03394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09133__A1 (.DIODE(_03394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09060__A1 (.DIODE(_03394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09669__B1 (.DIODE(_03395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09642__S1 (.DIODE(_03395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09623__B1 (.DIODE(_03395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09578__B1 (.DIODE(_03395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09529__S1 (.DIODE(_03395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09483__S1 (.DIODE(_03395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09303__S1 (.DIODE(_03395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09181__S1 (.DIODE(_03395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09130__S1 (.DIODE(_03395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09057__S1 (.DIODE(_03395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09646__S0 (.DIODE(_03400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09643__S0 (.DIODE(_03400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09533__S0 (.DIODE(_03400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09530__S0 (.DIODE(_03400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09487__S0 (.DIODE(_03400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09484__S0 (.DIODE(_03400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09307__S0 (.DIODE(_03400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09185__S0 (.DIODE(_03400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09134__S0 (.DIODE(_03400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09063__S0 (.DIODE(_03400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09646__S1 (.DIODE(_03401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09533__S1 (.DIODE(_03401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09487__S1 (.DIODE(_03401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09307__S1 (.DIODE(_03401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09186__S1 (.DIODE(_03401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09185__S1 (.DIODE(_03401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09135__S1 (.DIODE(_03401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09134__S1 (.DIODE(_03401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09064__S1 (.DIODE(_03401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09063__S1 (.DIODE(_03401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09469__A2 (.DIODE(_03408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09447__A2 (.DIODE(_03408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09402__A2 (.DIODE(_03408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09357__A2 (.DIODE(_03408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09335__A2 (.DIODE(_03408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09289__A2 (.DIODE(_03408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09244__A2 (.DIODE(_03408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09216__A2 (.DIODE(_03408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09167__A2 (.DIODE(_03408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09093__A2 (.DIODE(_03408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09707__S1 (.DIODE(_03418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09453__S1 (.DIODE(_03418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09431__S1 (.DIODE(_03418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09386__S1 (.DIODE(_03418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09345__S1 (.DIODE(_03418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09323__S1 (.DIODE(_03418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09277__S1 (.DIODE(_03418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09226__S1 (.DIODE(_03418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09202__S1 (.DIODE(_03418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09081__S1 (.DIODE(_03418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09092__B1 (.DIODE(_03429_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09093__C1 (.DIODE(_03430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09116__A2 (.DIODE(_03443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09139__A1 (.DIODE(_03474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09661__S0 (.DIODE(_03484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09615__S0 (.DIODE(_03484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09570__S0 (.DIODE(_03484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09548__S0 (.DIODE(_03484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09502__S0 (.DIODE(_03484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09456__S0 (.DIODE(_03484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09434__S0 (.DIODE(_03484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09389__S0 (.DIODE(_03484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09229__S0 (.DIODE(_03484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09151__S0 (.DIODE(_03484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09656__S1 (.DIODE(_03485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09615__S1 (.DIODE(_03485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09570__S1 (.DIODE(_03485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09548__S1 (.DIODE(_03485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09502__S1 (.DIODE(_03485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09456__S1 (.DIODE(_03485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09434__S1 (.DIODE(_03485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09389__S1 (.DIODE(_03485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09229__S1 (.DIODE(_03485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09151__S1 (.DIODE(_03485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09662__S0 (.DIODE(_03487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09616__S0 (.DIODE(_03487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09571__S0 (.DIODE(_03487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09549__S0 (.DIODE(_03487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09503__S0 (.DIODE(_03487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09457__S0 (.DIODE(_03487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09435__S0 (.DIODE(_03487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09390__S0 (.DIODE(_03487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09230__S0 (.DIODE(_03487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09154__S0 (.DIODE(_03487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09661__S1 (.DIODE(_03488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09616__S1 (.DIODE(_03488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09571__S1 (.DIODE(_03488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09549__S1 (.DIODE(_03488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09503__S1 (.DIODE(_03488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09457__S1 (.DIODE(_03488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09435__S1 (.DIODE(_03488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09390__S1 (.DIODE(_03488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09230__S1 (.DIODE(_03488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09154__S1 (.DIODE(_03488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09673__C1 (.DIODE(_03500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09627__C1 (.DIODE(_03500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09582__C1 (.DIODE(_03500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09560__C1 (.DIODE(_03500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09514__C1 (.DIODE(_03500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09468__C1 (.DIODE(_03500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09446__C1 (.DIODE(_03500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09401__C1 (.DIODE(_03500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09243__C1 (.DIODE(_03500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09166__C1 (.DIODE(_03500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09167__C1 (.DIODE(_03501_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09190__A1 (.DIODE(_03523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09707__S0 (.DIODE(_03534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09545__S0 (.DIODE(_03534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09453__S0 (.DIODE(_03534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09431__S0 (.DIODE(_03534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09386__S0 (.DIODE(_03534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09345__S0 (.DIODE(_03534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09323__S0 (.DIODE(_03534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09277__S0 (.DIODE(_03534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09226__S0 (.DIODE(_03534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09202__S0 (.DIODE(_03534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09711__S (.DIODE(_03539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09669__A1 (.DIODE(_03539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09623__A1 (.DIODE(_03539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09578__A1 (.DIODE(_03539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09556__A1 (.DIODE(_03539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09464__A1 (.DIODE(_03539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09442__A1 (.DIODE(_03539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09327__S (.DIODE(_03539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09281__S (.DIODE(_03539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09207__S (.DIODE(_03539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09715__A1 (.DIODE(_03543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09575__A1 (.DIODE(_03543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09553__A1 (.DIODE(_03543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09461__A1 (.DIODE(_03543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09439__A1 (.DIODE(_03543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09394__A1 (.DIODE(_03543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09331__A1 (.DIODE(_03543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09285__A1 (.DIODE(_03543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09235__A1 (.DIODE(_03543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09212__A1 (.DIODE(_03543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09216__C1 (.DIODE(_03548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09653__S0 (.DIODE(_03550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09607__S0 (.DIODE(_03550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09562__S0 (.DIODE(_03550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09540__S0 (.DIODE(_03550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09449__S0 (.DIODE(_03550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09448__S0 (.DIODE(_03550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09427__S0 (.DIODE(_03550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09426__S0 (.DIODE(_03550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09382__S0 (.DIODE(_03550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09220__S0 (.DIODE(_03550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09653__S1 (.DIODE(_03551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09607__S1 (.DIODE(_03551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09562__S1 (.DIODE(_03551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09540__S1 (.DIODE(_03551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09449__S1 (.DIODE(_03551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09448__S1 (.DIODE(_03551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09427__S1 (.DIODE(_03551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09426__S1 (.DIODE(_03551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09382__S1 (.DIODE(_03551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09220__S1 (.DIODE(_03551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09700__S0 (.DIODE(_03554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09656__S0 (.DIODE(_03554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09610__S0 (.DIODE(_03554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09565__S0 (.DIODE(_03554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09543__S0 (.DIODE(_03554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09496__S0 (.DIODE(_03554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09451__S0 (.DIODE(_03554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09429__S0 (.DIODE(_03554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09384__S0 (.DIODE(_03554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09224__S0 (.DIODE(_03554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09700__S1 (.DIODE(_03555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09610__S1 (.DIODE(_03555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09565__S1 (.DIODE(_03555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09543__S1 (.DIODE(_03555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09496__S1 (.DIODE(_03555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09451__S1 (.DIODE(_03555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09429__S1 (.DIODE(_03555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09384__S1 (.DIODE(_03555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09338__S1 (.DIODE(_03555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09224__S1 (.DIODE(_03555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09715__B1 (.DIODE(_03566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09666__B1 (.DIODE(_03566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09620__B1 (.DIODE(_03566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09575__B1 (.DIODE(_03566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09553__B1 (.DIODE(_03566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09461__B1 (.DIODE(_03566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09439__B1 (.DIODE(_03566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09394__B1 (.DIODE(_03566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09331__B1 (.DIODE(_03566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09235__B1 (.DIODE(_03566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09668__B_N (.DIODE(_03569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09622__B_N (.DIODE(_03569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09577__B_N (.DIODE(_03569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09555__B_N (.DIODE(_03569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09463__B_N (.DIODE(_03569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09441__B_N (.DIODE(_03569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09397__A1 (.DIODE(_03569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09396__B_N (.DIODE(_03569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09239__A1 (.DIODE(_03569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09238__B_N (.DIODE(_03569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09244__C1 (.DIODE(_03575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09267__B1 (.DIODE(_03597_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09271__A2 (.DIODE(_03600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09289__B2 (.DIODE(_03605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09312__A1 (.DIODE(_03640_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09317__A2 (.DIODE(_03644_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09335__B2 (.DIODE(_03649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09357__B2 (.DIODE(_03670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09380__B1 (.DIODE(_03705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09402__B2 (.DIODE(_03713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09447__B2 (.DIODE(_03756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09469__B2 (.DIODE(_03777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09538__A1 (.DIODE(_03856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09606__B1 (.DIODE(_03921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09651__A1 (.DIODE(_03964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09697__A3 (.DIODE(_04007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10768__S (.DIODE(_04034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10640__S (.DIODE(_04034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10593__S (.DIODE(_04034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10592__B (.DIODE(_04034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10591__A1 (.DIODE(_04034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10556__A2 (.DIODE(_04034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10555__A2 (.DIODE(_04034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10553__S (.DIODE(_04034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09756__A0 (.DIODE(_04034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09725__B1 (.DIODE(_04034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09872__C1 (.DIODE(_04041_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09754__A (.DIODE(_04041_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09735__A (.DIODE(_04041_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09855__C1 (.DIODE(_04042_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09843__C1 (.DIODE(_04042_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09838__C1 (.DIODE(_04042_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09826__C1 (.DIODE(_04042_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09795__C1 (.DIODE(_04042_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09790__C1 (.DIODE(_04042_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09785__C1 (.DIODE(_04042_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09767__C1 (.DIODE(_04042_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09749__B2 (.DIODE(_04042_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09736__B (.DIODE(_04042_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09737__A (.DIODE(_04043_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10273__B (.DIODE(_04045_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10232__B (.DIODE(_04045_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10228__B (.DIODE(_04045_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10182__A (.DIODE(_04045_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09893__B1 (.DIODE(_04045_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09861__A1 (.DIODE(_04045_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09860__A1 (.DIODE(_04045_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09831__A1 (.DIODE(_04045_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09741__A (.DIODE(_04045_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09893__C1 (.DIODE(_04046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09861__A2 (.DIODE(_04046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09860__A2 (.DIODE(_04046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09831__A2 (.DIODE(_04046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09741__B (.DIODE(_04046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09871__B (.DIODE(_04048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09854__B (.DIODE(_04048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09842__B (.DIODE(_04048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09837__B (.DIODE(_04048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09825__B (.DIODE(_04048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09794__B (.DIODE(_04048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09789__B (.DIODE(_04048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09784__B (.DIODE(_04048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09766__B (.DIODE(_04048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09743__A (.DIODE(_04048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09986__B1 (.DIODE(_04049_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09936__A (.DIODE(_04049_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09933__A (.DIODE(_04049_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09930__A (.DIODE(_04049_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09927__A (.DIODE(_04049_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09909__B1 (.DIODE(_04049_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09900__B1 (.DIODE(_04049_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09848__B1 (.DIODE(_04049_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09800__A2 (.DIODE(_04049_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09749__A1 (.DIODE(_04049_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09907__B (.DIODE(_04052_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09901__A (.DIODE(_04052_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09898__B (.DIODE(_04052_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09892__A1 (.DIODE(_04052_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09749__A2 (.DIODE(_04052_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09907__C (.DIODE(_04055_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09898__A_N (.DIODE(_04055_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09760__A3 (.DIODE(_04055_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09751__B (.DIODE(_04055_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09901__B_N (.DIODE(_04056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09892__A2 (.DIODE(_04056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09753__A1 (.DIODE(_04056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09938__A (.DIODE(_04057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09849__A (.DIODE(_04057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09832__A1 (.DIODE(_04057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09815__S (.DIODE(_04057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09810__S (.DIODE(_04057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09804__S (.DIODE(_04057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09777__A (.DIODE(_04057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09774__S (.DIODE(_04057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09765__B1 (.DIODE(_04057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09753__S (.DIODE(_04057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09888__S (.DIODE(_04059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09883__S (.DIODE(_04059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09878__S (.DIODE(_04059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09867__S (.DIODE(_04059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09862__S (.DIODE(_04059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09833__S (.DIODE(_04059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09816__S (.DIODE(_04059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09755__A (.DIODE(_04059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09873__A2 (.DIODE(_04060_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09856__A2 (.DIODE(_04060_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09850__B1 (.DIODE(_04060_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09821__B (.DIODE(_04060_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09811__S (.DIODE(_04060_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09805__S (.DIODE(_04060_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09800__C1 (.DIODE(_04060_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09775__S (.DIODE(_04060_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09758__A (.DIODE(_04060_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09756__S (.DIODE(_04060_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09757__A (.DIODE(_04061_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09851__A2_N (.DIODE(_04062_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09844__A2 (.DIODE(_04062_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09839__A2 (.DIODE(_04062_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09827__A2 (.DIODE(_04062_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09822__A1 (.DIODE(_04062_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09801__A2 (.DIODE(_04062_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09796__A2 (.DIODE(_04062_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09791__A2 (.DIODE(_04062_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09786__A2 (.DIODE(_04062_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09768__A2 (.DIODE(_04062_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09776__A (.DIODE(_04078_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09872__A1 (.DIODE(_04079_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09855__A1 (.DIODE(_04079_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09843__A1 (.DIODE(_04079_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09838__A1 (.DIODE(_04079_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09826__A1 (.DIODE(_04079_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09820__S (.DIODE(_04079_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09799__B1 (.DIODE(_04079_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09795__A1 (.DIODE(_04079_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09790__A1 (.DIODE(_04079_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09785__A1 (.DIODE(_04079_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10005__A (.DIODE(_04139_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10001__A (.DIODE(_04139_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09997__A (.DIODE(_04139_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09993__A (.DIODE(_04139_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09989__A (.DIODE(_04139_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09982__A (.DIODE(_04139_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09978__A (.DIODE(_04139_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09974__A (.DIODE(_04139_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09971__A (.DIODE(_04139_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09850__A2 (.DIODE(_04139_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09889__A (.DIODE(_04171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10591__B1 (.DIODE(_04173_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10192__A (.DIODE(_04173_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09984__B (.DIODE(_04173_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09902__A1 (.DIODE(_04173_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09895__A2 (.DIODE(_04173_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09892__B1 (.DIODE(_04173_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09902__B1 (.DIODE(_04175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09894__B (.DIODE(_04175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09948__A2 (.DIODE(_04176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09945__A2 (.DIODE(_04176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09942__A2 (.DIODE(_04176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09939__A2 (.DIODE(_04176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09935__A2 (.DIODE(_04176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09932__A2 (.DIODE(_04176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09929__A2 (.DIODE(_04176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09926__A2 (.DIODE(_04176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09900__A1 (.DIODE(_04176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11374__C1 (.DIODE(_04177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11308__C1 (.DIODE(_04177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11251__C1 (.DIODE(_04177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11178__B1 (.DIODE(_04177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11088__C1 (.DIODE(_04177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11041__C1 (.DIODE(_04177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10974__C1 (.DIODE(_04177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10885__C1 (.DIODE(_04177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10547__A (.DIODE(_04177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09897__A (.DIODE(_04177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11646__B1 (.DIODE(_04178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11539__C1 (.DIODE(_04178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11517__A (.DIODE(_04178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11496__C1 (.DIODE(_04178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11474__A1 (.DIODE(_04178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11423__C1 (.DIODE(_04178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11347__A (.DIODE(_04178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11278__B1 (.DIODE(_04178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09907__A (.DIODE(_04178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09898__C (.DIODE(_04178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09948__B1 (.DIODE(_04180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09945__B1 (.DIODE(_04180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09942__B1 (.DIODE(_04180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09939__B1 (.DIODE(_04180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09935__B1 (.DIODE(_04180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09932__B1 (.DIODE(_04180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09929__B1 (.DIODE(_04180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09926__B1 (.DIODE(_04180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09900__A2 (.DIODE(_04180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11438__A2 (.DIODE(_04183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11407__A2 (.DIODE(_04183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11164__A2 (.DIODE(_04183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10003__A2 (.DIODE(_04183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09999__A2 (.DIODE(_04183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09995__A2 (.DIODE(_04183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09991__A2 (.DIODE(_04183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09987__A2 (.DIODE(_04183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09980__A2 (.DIODE(_04183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09905__A (.DIODE(_04183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09976__A2 (.DIODE(_04184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09973__A2 (.DIODE(_04184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09970__A2 (.DIODE(_04184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09967__A2 (.DIODE(_04184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09964__A2 (.DIODE(_04184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09961__A2 (.DIODE(_04184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09958__A2 (.DIODE(_04184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09955__A2 (.DIODE(_04184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09952__A2 (.DIODE(_04184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09909__A1 (.DIODE(_04184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09968__A (.DIODE(_04204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09965__A (.DIODE(_04204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09962__A (.DIODE(_04204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09959__A (.DIODE(_04204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09956__A (.DIODE(_04204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09953__A (.DIODE(_04204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09949__A (.DIODE(_04204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09946__A (.DIODE(_04204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09943__A (.DIODE(_04204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09940__A (.DIODE(_04204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09973__B1 (.DIODE(_04213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09970__B1 (.DIODE(_04213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09967__B1 (.DIODE(_04213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09964__B1 (.DIODE(_04213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09961__B1 (.DIODE(_04213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09958__B1 (.DIODE(_04213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09955__B1 (.DIODE(_04213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09952__B1 (.DIODE(_04213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10273__C (.DIODE(_04360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10232__C (.DIODE(_04360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10228__C (.DIODE(_04360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10182__B (.DIODE(_04360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10179__B (.DIODE(_04360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11121__A2 (.DIODE(_04361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11057__A (.DIODE(_04361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10186__A (.DIODE(_04361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10687__A (.DIODE(_04363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10615__S (.DIODE(_04363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10599__A (.DIODE(_04363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10546__A (.DIODE(_04363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10545__B1 (.DIODE(_04363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10538__S (.DIODE(_04363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10466__S (.DIODE(_04363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10463__S (.DIODE(_04363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10438__S (.DIODE(_04363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10184__A (.DIODE(_04363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10288__S (.DIODE(_04364_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10262__S (.DIODE(_04364_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10245__S (.DIODE(_04364_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10236__S (.DIODE(_04364_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10221__S (.DIODE(_04364_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10183__A (.DIODE(_04364_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11215__A1 (.DIODE(_04365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10728__S (.DIODE(_04365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10546__B (.DIODE(_04365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10545__A1 (.DIODE(_04365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10303__S (.DIODE(_04365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10298__S (.DIODE(_04365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10290__S (.DIODE(_04365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10253__S (.DIODE(_04365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10224__S (.DIODE(_04365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10184__B (.DIODE(_04365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11474__A2 (.DIODE(_04366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11347__B (.DIODE(_04366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11227__A1 (.DIODE(_04366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10673__B (.DIODE(_04366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10600__A (.DIODE(_04366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10186__B (.DIODE(_04366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11365__B1 (.DIODE(_04375_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11329__B1 (.DIODE(_04375_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11296__B1 (.DIODE(_04375_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11241__B1 (.DIODE(_04375_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11224__B1 (.DIODE(_04375_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11136__B1 (.DIODE(_04375_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10850__B1 (.DIODE(_04375_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10811__B1 (.DIODE(_04375_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10721__B1 (.DIODE(_04375_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10194__A (.DIODE(_04375_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11604__B1 (.DIODE(_04376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11547__B1 (.DIODE(_04376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11436__A1 (.DIODE(_04376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11188__B1 (.DIODE(_04376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11010__B1 (.DIODE(_04376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10980__B1 (.DIODE(_04376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10901__B2 (.DIODE(_04376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10675__A1 (.DIODE(_04376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10633__B1 (.DIODE(_04376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10550__A1 (.DIODE(_04376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11364__A2 (.DIODE(_04384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11323__A2 (.DIODE(_04384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11295__A2 (.DIODE(_04384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11240__A2 (.DIODE(_04384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11223__A2 (.DIODE(_04384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11134__A2 (.DIODE(_04384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10849__A2 (.DIODE(_04384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10810__A2 (.DIODE(_04384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10596__A2 (.DIODE(_04384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10203__A (.DIODE(_04384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11651__A2 (.DIODE(_04385_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11603__A2 (.DIODE(_04385_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11546__A2 (.DIODE(_04385_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11434__A2 (.DIODE(_04385_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11187__A2 (.DIODE(_04385_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11009__A2 (.DIODE(_04385_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10979__A2 (.DIODE(_04385_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10900__A2 (.DIODE(_04385_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10644__A2 (.DIODE(_04385_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10218__A2 (.DIODE(_04385_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11469__B1 (.DIODE(_04388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11119__B1 (.DIODE(_04388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11058__A2 (.DIODE(_04388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10761__A (.DIODE(_04388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10207__A (.DIODE(_04388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11363__B1 (.DIODE(_04389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11322__B1 (.DIODE(_04389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11294__B1 (.DIODE(_04389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11239__B1 (.DIODE(_04389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11222__B1 (.DIODE(_04389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11133__A2 (.DIODE(_04389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10848__B1 (.DIODE(_04389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10809__A2 (.DIODE(_04389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10719__A2 (.DIODE(_04389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10208__A (.DIODE(_04389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11650__B1 (.DIODE(_04390_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11602__B1 (.DIODE(_04390_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11545__B1 (.DIODE(_04390_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11433__B1 (.DIODE(_04390_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11186__B1 (.DIODE(_04390_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10978__B1 (.DIODE(_04390_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10899__B1 (.DIODE(_04390_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10643__A2 (.DIODE(_04390_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10597__B1 (.DIODE(_04390_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10218__B1 (.DIODE(_04390_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11469__A2 (.DIODE(_04391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11322__A2 (.DIODE(_04391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11222__A2 (.DIODE(_04391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11119__A2 (.DIODE(_04391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10210__A (.DIODE(_04391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11390__A2 (.DIODE(_04392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11363__A2 (.DIODE(_04392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11294__A2 (.DIODE(_04392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11263__A2 (.DIODE(_04392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11239__A2 (.DIODE(_04392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11059__B1 (.DIODE(_04392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10941__A2 (.DIODE(_04392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10898__A (.DIODE(_04392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10848__A2 (.DIODE(_04392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10211__A (.DIODE(_04392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11602__A2 (.DIODE(_04393_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11545__A2 (.DIODE(_04393_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11433__A2 (.DIODE(_04393_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11009__B1 (.DIODE(_04393_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10810__B1 (.DIODE(_04393_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10763__B1 (.DIODE(_04393_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10720__B1 (.DIODE(_04393_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10644__B1 (.DIODE(_04393_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10597__A2 (.DIODE(_04393_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10217__A2 (.DIODE(_04393_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11627__B1 (.DIODE(_04395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11484__B1 (.DIODE(_04395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11391__B1 (.DIODE(_04395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11264__B1 (.DIODE(_04395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11240__B1 (.DIODE(_04395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10942__B1 (.DIODE(_04395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10849__B1 (.DIODE(_04395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10643__B1 (.DIODE(_04395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10596__B1 (.DIODE(_04395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10217__B1 (.DIODE(_04395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10217__C1 (.DIODE(_04398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11282__C1 (.DIODE(_04401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11116__C1 (.DIODE(_04401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11089__A1 (.DIODE(_04401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10714__C1 (.DIODE(_04401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10673__A (.DIODE(_04401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10630__C1 (.DIODE(_04401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10220__A (.DIODE(_04401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11625__A (.DIODE(_04402_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11576__A1_N (.DIODE(_04402_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11405__A1 (.DIODE(_04402_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11220__A (.DIODE(_04402_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11216__C1 (.DIODE(_04402_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11157__A1 (.DIODE(_04402_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11007__A1_N (.DIODE(_04402_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10940__A1_N (.DIODE(_04402_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10847__A1_N (.DIODE(_04402_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10549__A1 (.DIODE(_04402_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10269__A2 (.DIODE(_04408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10268__B (.DIODE(_04408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10231__A2 (.DIODE(_04408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10227__A2 (.DIODE(_04408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10278__A (.DIODE(_04450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10270__A2 (.DIODE(_04450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10272__A (.DIODE(_04451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10270__B1 (.DIODE(_04451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11003__B1 (.DIODE(_04480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10955__A2 (.DIODE(_04480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10309__A2 (.DIODE(_04480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10300__B (.DIODE(_04480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10299__B (.DIODE(_04480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11003__A2 (.DIODE(_04485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10973__B (.DIODE(_04485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10972__B (.DIODE(_04485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10305__B (.DIODE(_04485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10304__B (.DIODE(_04485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11584__B1 (.DIODE(_04498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10411__B1 (.DIODE(_04498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10409__B1 (.DIODE(_04498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10405__B1 (.DIODE(_04498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10402__B1 (.DIODE(_04498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10398__B1 (.DIODE(_04498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10382__B1 (.DIODE(_04498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10341__B1 (.DIODE(_04498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10339__B1 (.DIODE(_04498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10317__A (.DIODE(_04498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11584__A2 (.DIODE(_04520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11085__A1 (.DIODE(_04520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10670__A (.DIODE(_04520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10606__A (.DIODE(_04520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10411__A2 (.DIODE(_04520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10409__A2 (.DIODE(_04520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10405__A2 (.DIODE(_04520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10398__A2 (.DIODE(_04520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10382__A2 (.DIODE(_04520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10339__A2 (.DIODE(_04520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11452__B1 (.DIODE(_04547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10432__B (.DIODE(_04547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10366__B1 (.DIODE(_04547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10416__A2 (.DIODE(_04559_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10608__B (.DIODE(_04617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10605__B (.DIODE(_04617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10598__B (.DIODE(_04617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10545__A2 (.DIODE(_04617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10436__B (.DIODE(_04617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11138__S (.DIODE(_04620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11070__S (.DIODE(_04620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10526__A (.DIODE(_04620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10439__A (.DIODE(_04620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10531__A (.DIODE(_04626_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10510__S (.DIODE(_04626_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10492__A (.DIODE(_04626_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10489__S (.DIODE(_04626_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10474__S (.DIODE(_04626_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10457__S (.DIODE(_04626_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10445__A (.DIODE(_04626_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10911__A (.DIODE(_04633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10875__S (.DIODE(_04633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10795__S (.DIODE(_04633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10750__S (.DIODE(_04633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10530__A (.DIODE(_04633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10452__A (.DIODE(_04633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11063__S (.DIODE(_04645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11031__S (.DIODE(_04645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10987__S (.DIODE(_04645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10965__S (.DIODE(_04645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10958__A (.DIODE(_04645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10912__A1 (.DIODE(_04645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10829__A1 (.DIODE(_04645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10464__A (.DIODE(_04645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11032__C1 (.DIODE(_04648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10877__S (.DIODE(_04648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10797__S (.DIODE(_04648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10504__A (.DIODE(_04648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10483__A (.DIODE(_04648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10467__A (.DIODE(_04648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10911__B (.DIODE(_04659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10533__A (.DIODE(_04659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10529__B (.DIODE(_04659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10478__A1 (.DIODE(_04659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11622__A0 (.DIODE(_04723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11561__A1 (.DIODE(_04723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11515__A0 (.DIODE(_04723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11394__A0 (.DIODE(_04723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11318__A0 (.DIODE(_04723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11217__A0 (.DIODE(_04723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10998__A0 (.DIODE(_04723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10756__A0 (.DIODE(_04723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10649__A0 (.DIODE(_04723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10543__A1 (.DIODE(_04723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11403__B1 (.DIODE(_04729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11376__A1 (.DIODE(_04729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11099__B1 (.DIODE(_04729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10931__B1 (.DIODE(_04729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10896__C1 (.DIODE(_04729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10843__B1 (.DIODE(_04729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10808__A1 (.DIODE(_04729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10685__A (.DIODE(_04729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10607__B1 (.DIODE(_04729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10548__B1 (.DIODE(_04729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10550__B1_N (.DIODE(_04731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10864__A1 (.DIODE(_04734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10819__A (.DIODE(_04734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10778__A (.DIODE(_04734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10769__A (.DIODE(_04734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10682__A (.DIODE(_04734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10641__A (.DIODE(_04734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10594__A (.DIODE(_04734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10557__B1 (.DIODE(_04734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10592__A_N (.DIODE(_04736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10591__A2 (.DIODE(_04736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10555__B1 (.DIODE(_04736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11633__A1 (.DIODE(_04741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11579__A1 (.DIODE(_04741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11526__A1 (.DIODE(_04741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11501__A1 (.DIODE(_04741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11476__A1 (.DIODE(_04741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11349__A1 (.DIODE(_04741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11286__A1 (.DIODE(_04741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10767__A (.DIODE(_04741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10563__B (.DIODE(_04741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10560__B (.DIODE(_04741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10572__A4 (.DIODE(_04753_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14114__A (.DIODE(_04755_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14103__A (.DIODE(_04755_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14024__A (.DIODE(_04755_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14013__A (.DIODE(_04755_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14002__A (.DIODE(_04755_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13891__A (.DIODE(_04755_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12112__A (.DIODE(_04755_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12110__A (.DIODE(_04755_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10574__B1 (.DIODE(_04755_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11765__B (.DIODE(_04756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10583__A (.DIODE(_04756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10581__B (.DIODE(_04756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10577__A1 (.DIODE(_04756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10576__B1 (.DIODE(_04756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11634__A (.DIODE(_04759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11580__A (.DIODE(_04759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11527__A (.DIODE(_04759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11502__A (.DIODE(_04759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11477__A (.DIODE(_04759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11287__A (.DIODE(_04759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11233__A (.DIODE(_04759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10590__A (.DIODE(_04759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10578__A (.DIODE(_04759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14035__A1 (.DIODE(_04761_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12529__A (.DIODE(_04761_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11663__A (.DIODE(_04761_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10580__A (.DIODE(_04761_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13516__A0 (.DIODE(_04762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13380__A0 (.DIODE(_04762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13312__A0 (.DIODE(_04762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13244__A0 (.DIODE(_04762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12971__A0 (.DIODE(_04762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12699__A0 (.DIODE(_04762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12326__A0 (.DIODE(_04762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12044__A0 (.DIODE(_04762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11769__A0 (.DIODE(_04762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10588__A0 (.DIODE(_04762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11661__S (.DIODE(_04768_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11636__S (.DIODE(_04768_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11353__A (.DIODE(_04768_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11016__A (.DIODE(_04768_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10587__A (.DIODE(_04768_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10985__S (.DIODE(_04769_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10948__S (.DIODE(_04769_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10906__S (.DIODE(_04769_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10855__S (.DIODE(_04769_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10816__S (.DIODE(_04769_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10775__S (.DIODE(_04769_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10726__S (.DIODE(_04769_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10679__S (.DIODE(_04769_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10638__S (.DIODE(_04769_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10588__S (.DIODE(_04769_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11659__C1 (.DIODE(_04771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11440__C1 (.DIODE(_04771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11409__C1 (.DIODE(_04771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11092__A (.DIODE(_04771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10946__A (.DIODE(_04771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10853__A (.DIODE(_04771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10814__A (.DIODE(_04771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10724__A (.DIODE(_04771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10677__A (.DIODE(_04771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10636__A (.DIODE(_04771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11641__B1 (.DIODE(_04782_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11621__A1 (.DIODE(_04782_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11512__A1 (.DIODE(_04782_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11489__A (.DIODE(_04782_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11399__B1 (.DIODE(_04782_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11244__A (.DIODE(_04782_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10953__B (.DIODE(_04782_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10738__A1 (.DIODE(_04782_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10672__A1 (.DIODE(_04782_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10602__B1 (.DIODE(_04782_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11345__A (.DIODE(_04786_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11274__A1 (.DIODE(_04786_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11214__A (.DIODE(_04786_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11085__B1 (.DIODE(_04786_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10670__B (.DIODE(_04786_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10606__B (.DIODE(_04786_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11303__B2 (.DIODE(_04787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11246__B1 (.DIODE(_04787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11101__B1 (.DIODE(_04787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10931__A1 (.DIODE(_04787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10895__A (.DIODE(_04787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10843__A1 (.DIODE(_04787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10607__A3 (.DIODE(_04787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11466__A1 (.DIODE(_04808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11145__A1 (.DIODE(_04808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11116__A1 (.DIODE(_04808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11073__A1 (.DIODE(_04808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10925__A1 (.DIODE(_04808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10836__A1 (.DIODE(_04808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10647__A (.DIODE(_04808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10628__A1 (.DIODE(_04808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10633__C1 (.DIODE(_04813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11633__B1 (.DIODE(_04815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11579__B1 (.DIODE(_04815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11312__B2 (.DIODE(_04815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11257__B2 (.DIODE(_04815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11159__B2 (.DIODE(_04815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11125__B2 (.DIODE(_04815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11091__B2 (.DIODE(_04815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10723__B2 (.DIODE(_04815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10676__B2 (.DIODE(_04815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10635__B2 (.DIODE(_04815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14037__A1 (.DIODE(_04817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12534__A (.DIODE(_04817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11670__A (.DIODE(_04817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10637__A (.DIODE(_04817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13518__A0 (.DIODE(_04818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13382__A0 (.DIODE(_04818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13314__A0 (.DIODE(_04818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13246__A0 (.DIODE(_04818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12973__A0 (.DIODE(_04818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12701__A0 (.DIODE(_04818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12328__A0 (.DIODE(_04818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12046__A0 (.DIODE(_04818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11771__A0 (.DIODE(_04818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10638__A0 (.DIODE(_04818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11628__B1 (.DIODE(_04825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11522__C (.DIODE(_04825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11267__B1 (.DIODE(_04825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11131__A (.DIODE(_04825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11122__A3 (.DIODE(_04825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11048__A2 (.DIODE(_04825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10980__A2 (.DIODE(_04825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10765__A2 (.DIODE(_04825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10684__A (.DIODE(_04825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10646__A1 (.DIODE(_04825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11622__A1 (.DIODE(_04827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11588__A1 (.DIODE(_04827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11561__A0 (.DIODE(_04827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11515__A1 (.DIODE(_04827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11394__A1 (.DIODE(_04827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11318__A1 (.DIODE(_04827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11217__A1 (.DIODE(_04827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10998__A1 (.DIODE(_04827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10756__A1 (.DIODE(_04827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10649__A1 (.DIODE(_04827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11497__A1 (.DIODE(_04831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11424__A1 (.DIODE(_04831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11375__A1 (.DIODE(_04831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11309__A1 (.DIODE(_04831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11252__A1 (.DIODE(_04831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11179__B2 (.DIODE(_04831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11042__A1 (.DIODE(_04831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10975__A1 (.DIODE(_04831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10886__A1 (.DIODE(_04831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10652__B (.DIODE(_04831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11429__B1 (.DIODE(_04850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10782__B1 (.DIODE(_04850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10691__A (.DIODE(_04850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10671__B1 (.DIODE(_04850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11620__B1 (.DIODE(_04853_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11542__A1 (.DIODE(_04853_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11511__B1 (.DIODE(_04853_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11472__A1 (.DIODE(_04853_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11430__B1 (.DIODE(_04853_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11254__A1 (.DIODE(_04853_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11156__C1 (.DIODE(_04853_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10977__A1 (.DIODE(_04853_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10759__A1 (.DIODE(_04853_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10674__B2 (.DIODE(_04853_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10675__C1 (.DIODE(_04854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14039__A1 (.DIODE(_04857_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12537__A (.DIODE(_04857_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11673__A (.DIODE(_04857_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10678__A (.DIODE(_04857_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13520__A0 (.DIODE(_04858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13384__A0 (.DIODE(_04858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13316__A0 (.DIODE(_04858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13248__A0 (.DIODE(_04858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12975__A0 (.DIODE(_04858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12703__A0 (.DIODE(_04858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12330__A0 (.DIODE(_04858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12048__A0 (.DIODE(_04858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11773__A0 (.DIODE(_04858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10679__A0 (.DIODE(_04858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11465__B1 (.DIODE(_04863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11377__A1 (.DIODE(_04863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11311__A1 (.DIODE(_04863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11226__A1 (.DIODE(_04863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11010__A2 (.DIODE(_04863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10944__A2 (.DIODE(_04863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10867__B (.DIODE(_04863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10851__A2 (.DIODE(_04863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10812__A2 (.DIODE(_04863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10722__A2 (.DIODE(_04863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11656__A1 (.DIODE(_04864_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11598__B2 (.DIODE(_04864_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11576__B1 (.DIODE(_04864_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11498__A1 (.DIODE(_04864_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11321__B1 (.DIODE(_04864_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11310__A1 (.DIODE(_04864_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11182__A1 (.DIODE(_04864_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11025__C1 (.DIODE(_04864_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11007__B1 (.DIODE(_04864_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10716__A1 (.DIODE(_04864_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11367__C1 (.DIODE(_04867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11303__A1 (.DIODE(_04867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11099__A1 (.DIODE(_04867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10939__C (.DIODE(_04867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10891__B1 (.DIODE(_04867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10689__A (.DIODE(_04867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11597__B2 (.DIODE(_04868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11575__A1 (.DIODE(_04868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11533__B1 (.DIODE(_04868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11431__A1 (.DIODE(_04868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11171__A1 (.DIODE(_04868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11024__A (.DIODE(_04868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11002__B1 (.DIODE(_04868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10846__C1 (.DIODE(_04868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10786__C1 (.DIODE(_04868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10690__C1 (.DIODE(_04868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11645__A (.DIODE(_04870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11619__B1 (.DIODE(_04870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11536__B2 (.DIODE(_04870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11511__A1 (.DIODE(_04870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11371__B1 (.DIODE(_04870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11278__A1 (.DIODE(_04870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11169__B1 (.DIODE(_04870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11156__A1 (.DIODE(_04870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10737__B1 (.DIODE(_04870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10692__B1 (.DIODE(_04870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11175__B1 (.DIODE(_04879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11173__B1 (.DIODE(_04879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11143__B1 (.DIODE(_04879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11071__B1 (.DIODE(_04879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11036__B1 (.DIODE(_04879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10861__A (.DIODE(_04879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10833__B1 (.DIODE(_04879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10800__B1 (.DIODE(_04879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10745__B1 (.DIODE(_04879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10701__C1 (.DIODE(_04879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11539__A1 (.DIODE(_04891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11496__A1 (.DIODE(_04891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11423__B2 (.DIODE(_04891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11374__A1 (.DIODE(_04891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11308__B2 (.DIODE(_04891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11178__A2 (.DIODE(_04891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11041__B2 (.DIODE(_04891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10974__B2 (.DIODE(_04891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10885__B2 (.DIODE(_04891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10713__A (.DIODE(_04891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10722__B1 (.DIODE(_04895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11627__A2 (.DIODE(_04896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11558__A2 (.DIODE(_04896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11519__A2 (.DIODE(_04896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11484__A2 (.DIODE(_04896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11391__A2 (.DIODE(_04896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11264__A2 (.DIODE(_04896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11046__A2 (.DIODE(_04896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10942__A2 (.DIODE(_04896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10763__A2 (.DIODE(_04896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10720__A2 (.DIODE(_04896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11470__B1 (.DIODE(_04897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11364__B1 (.DIODE(_04897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11323__B1 (.DIODE(_04897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11295__B1 (.DIODE(_04897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11223__B1 (.DIODE(_04897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11008__B1 (.DIODE(_04897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10897__A (.DIODE(_04897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10809__B1 (.DIODE(_04897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10762__B1 (.DIODE(_04897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10719__B1 (.DIODE(_04897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14041__A1 (.DIODE(_04903_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12540__A (.DIODE(_04903_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11676__A (.DIODE(_04903_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10725__A (.DIODE(_04903_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13522__A0 (.DIODE(_04904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13386__A0 (.DIODE(_04904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13318__A0 (.DIODE(_04904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13250__A0 (.DIODE(_04904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12977__A0 (.DIODE(_04904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12705__A0 (.DIODE(_04904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12332__A0 (.DIODE(_04904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12050__A0 (.DIODE(_04904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11775__A0 (.DIODE(_04904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10726__A0 (.DIODE(_04904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11624__A1 (.DIODE(_04917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11564__B2 (.DIODE(_04917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11513__A (.DIODE(_04917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11396__A1 (.DIODE(_04917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11317__A (.DIODE(_04917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11219__B2 (.DIODE(_04917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11136__A1 (.DIODE(_04917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11000__A1 (.DIODE(_04917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10888__A1 (.DIODE(_04917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10758__A1 (.DIODE(_04917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11626__B1 (.DIODE(_04939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11557__B1 (.DIODE(_04939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11518__B1 (.DIODE(_04939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11483__B1 (.DIODE(_04939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11390__B1 (.DIODE(_04939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11263__B1 (.DIODE(_04939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11045__B1 (.DIODE(_04939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11008__A2 (.DIODE(_04939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10941__B1 (.DIODE(_04939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10762__A2 (.DIODE(_04939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14043__A1 (.DIODE(_04951_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12543__A (.DIODE(_04951_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11679__A (.DIODE(_04951_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10774__A (.DIODE(_04951_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13524__A0 (.DIODE(_04952_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13388__A0 (.DIODE(_04952_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13320__A0 (.DIODE(_04952_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13252__A0 (.DIODE(_04952_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12979__A0 (.DIODE(_04952_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12707__A0 (.DIODE(_04952_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12334__A0 (.DIODE(_04952_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12052__A0 (.DIODE(_04952_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11777__A0 (.DIODE(_04952_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10775__A0 (.DIODE(_04952_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10812__B1 (.DIODE(_04985_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10811__B2 (.DIODE(_04987_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14045__A1 (.DIODE(_04991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12546__A (.DIODE(_04991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11682__A (.DIODE(_04991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10815__A (.DIODE(_04991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13526__A0 (.DIODE(_04992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13390__A0 (.DIODE(_04992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13322__A0 (.DIODE(_04992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13254__A0 (.DIODE(_04992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12981__A0 (.DIODE(_04992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12709__A0 (.DIODE(_04992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12336__A0 (.DIODE(_04992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12054__A0 (.DIODE(_04992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11779__A0 (.DIODE(_04992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10816__A0 (.DIODE(_04992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10851__B1 (.DIODE(_05023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14047__A1 (.DIODE(_05029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12549__A (.DIODE(_05029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11685__A (.DIODE(_05029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10854__A (.DIODE(_05029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13528__A0 (.DIODE(_05030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13392__A0 (.DIODE(_05030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13324__A0 (.DIODE(_05030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13256__A0 (.DIODE(_05030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12983__A0 (.DIODE(_05030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12711__A0 (.DIODE(_05030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12338__A0 (.DIODE(_05030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12056__A0 (.DIODE(_05030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11781__A0 (.DIODE(_05030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10855__A0 (.DIODE(_05030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11608__A (.DIODE(_05032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11551__A (.DIODE(_05032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11191__A (.DIODE(_05032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10983__A (.DIODE(_05032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10904__A (.DIODE(_05032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11539__B2 (.DIODE(_05057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11496__B2 (.DIODE(_05057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11423__A1 (.DIODE(_05057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11374__B2 (.DIODE(_05057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11308__A1 (.DIODE(_05057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11251__B2 (.DIODE(_05057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11179__A1 (.DIODE(_05057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11041__A1 (.DIODE(_05057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10974__A1 (.DIODE(_05057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10885__A1 (.DIODE(_05057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10901__A1 (.DIODE(_05063_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11597__A1 (.DIODE(_05070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11575__B2 (.DIODE(_05070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11493__B2 (.DIODE(_05070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11459__A (.DIODE(_05070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11403__A1 (.DIODE(_05070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11344__B1 (.DIODE(_05070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11025__A1 (.DIODE(_05070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11006__B2 (.DIODE(_05070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10956__B1 (.DIODE(_05070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10896__B2 (.DIODE(_05070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10901__A2 (.DIODE(_05071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11650__A2 (.DIODE(_05073_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11626__A2 (.DIODE(_05073_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11557__A2 (.DIODE(_05073_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11518__A2 (.DIODE(_05073_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11483__A2 (.DIODE(_05073_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11186__A2 (.DIODE(_05073_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11134__B1 (.DIODE(_05073_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11045__A2 (.DIODE(_05073_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10978__A2 (.DIODE(_05073_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10899__A2 (.DIODE(_05073_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10901__B1 (.DIODE(_05075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14049__A1 (.DIODE(_05079_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12552__A (.DIODE(_05079_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11688__A (.DIODE(_05079_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10905__A (.DIODE(_05079_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13530__A0 (.DIODE(_05080_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13394__A0 (.DIODE(_05080_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13326__A0 (.DIODE(_05080_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13258__A0 (.DIODE(_05080_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12985__A0 (.DIODE(_05080_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12713__A0 (.DIODE(_05080_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12340__A0 (.DIODE(_05080_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12058__A0 (.DIODE(_05080_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11783__A0 (.DIODE(_05080_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10906__A0 (.DIODE(_05080_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10944__B1 (.DIODE(_05114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14051__A1 (.DIODE(_05120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12555__A (.DIODE(_05120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11691__A (.DIODE(_05120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10947__A (.DIODE(_05120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13532__A0 (.DIODE(_05121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13396__A0 (.DIODE(_05121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13328__A0 (.DIODE(_05121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13260__A0 (.DIODE(_05121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12987__A0 (.DIODE(_05121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12715__A0 (.DIODE(_05121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12342__A0 (.DIODE(_05121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12060__A0 (.DIODE(_05121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11785__A0 (.DIODE(_05121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10948__A0 (.DIODE(_05121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10981__B1 (.DIODE(_05150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10980__B2 (.DIODE(_05152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14053__A1 (.DIODE(_05156_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12558__A (.DIODE(_05156_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11694__A (.DIODE(_05156_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10984__A (.DIODE(_05156_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13534__A0 (.DIODE(_05157_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13398__A0 (.DIODE(_05157_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13330__A0 (.DIODE(_05157_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13262__A0 (.DIODE(_05157_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12989__A0 (.DIODE(_05157_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12717__A0 (.DIODE(_05157_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12344__A0 (.DIODE(_05157_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12062__A0 (.DIODE(_05157_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11787__A0 (.DIODE(_05157_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10985__A0 (.DIODE(_05157_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11011__B1 (.DIODE(_05179_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14056__A1 (.DIODE(_05186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12561__A (.DIODE(_05186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11697__A (.DIODE(_05186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11015__A (.DIODE(_05186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13537__A0 (.DIODE(_05187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13401__A0 (.DIODE(_05187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13333__A0 (.DIODE(_05187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13265__A0 (.DIODE(_05187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12992__A0 (.DIODE(_05187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12720__A0 (.DIODE(_05187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12347__A0 (.DIODE(_05187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12065__A0 (.DIODE(_05187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11790__A0 (.DIODE(_05187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11017__A0 (.DIODE(_05187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11315__S (.DIODE(_05188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11289__S (.DIODE(_05188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11260__S (.DIODE(_05188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11235__S (.DIODE(_05188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11193__S (.DIODE(_05188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11162__S (.DIODE(_05188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11128__S (.DIODE(_05188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11094__S (.DIODE(_05188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11054__S (.DIODE(_05188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11017__S (.DIODE(_05188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11049__A1 (.DIODE(_05196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11048__B2 (.DIODE(_05217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14058__A1 (.DIODE(_05223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12565__A (.DIODE(_05223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11701__A (.DIODE(_05223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11053__A (.DIODE(_05223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13539__A0 (.DIODE(_05224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13403__A0 (.DIODE(_05224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13335__A0 (.DIODE(_05224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13267__A0 (.DIODE(_05224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12994__A0 (.DIODE(_05224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12722__A0 (.DIODE(_05224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12349__A0 (.DIODE(_05224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12067__A0 (.DIODE(_05224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11792__A0 (.DIODE(_05224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11054__A0 (.DIODE(_05224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11061__B2 (.DIODE(_05229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11090__C_N (.DIODE(_05259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14060__A1 (.DIODE(_05262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12568__A (.DIODE(_05262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11704__A (.DIODE(_05262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11093__A (.DIODE(_05262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13541__A0 (.DIODE(_05263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13405__A0 (.DIODE(_05263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13337__A0 (.DIODE(_05263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13269__A0 (.DIODE(_05263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12996__A0 (.DIODE(_05263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12724__A0 (.DIODE(_05263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12351__A0 (.DIODE(_05263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12069__A0 (.DIODE(_05263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11794__A0 (.DIODE(_05263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11094__A0 (.DIODE(_05263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11124__A (.DIODE(_05287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11121__B2 (.DIODE(_05289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14062__A1 (.DIODE(_05295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12571__A (.DIODE(_05295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11707__A (.DIODE(_05295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11127__A (.DIODE(_05295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13543__A0 (.DIODE(_05296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13407__A0 (.DIODE(_05296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13339__A0 (.DIODE(_05296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13271__A0 (.DIODE(_05296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12998__A0 (.DIODE(_05296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12726__A0 (.DIODE(_05296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12353__A0 (.DIODE(_05296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12071__A0 (.DIODE(_05296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11796__A0 (.DIODE(_05296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11128__A0 (.DIODE(_05296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11136__B2 (.DIODE(_05302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11158__C1 (.DIODE(_05325_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14064__A1 (.DIODE(_05328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12574__A (.DIODE(_05328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11710__A (.DIODE(_05328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11161__A (.DIODE(_05328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13545__A0 (.DIODE(_05329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13409__A0 (.DIODE(_05329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13341__A0 (.DIODE(_05329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13273__A0 (.DIODE(_05329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13000__A0 (.DIODE(_05329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12728__A0 (.DIODE(_05329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12355__A0 (.DIODE(_05329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12073__A0 (.DIODE(_05329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11798__A0 (.DIODE(_05329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11162__A0 (.DIODE(_05329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11190__B1 (.DIODE(_05349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11188__B2 (.DIODE(_05354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14066__A1 (.DIODE(_05358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12577__A (.DIODE(_05358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11713__A (.DIODE(_05358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11192__A (.DIODE(_05358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13547__A0 (.DIODE(_05359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13411__A0 (.DIODE(_05359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13343__A0 (.DIODE(_05359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13275__A0 (.DIODE(_05359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13002__A0 (.DIODE(_05359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12730__A0 (.DIODE(_05359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12357__A0 (.DIODE(_05359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12075__A0 (.DIODE(_05359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11800__A0 (.DIODE(_05359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11193__A0 (.DIODE(_05359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11227__A2 (.DIODE(_05382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11224__B2 (.DIODE(_05389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14068__A1 (.DIODE(_05399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12580__A (.DIODE(_05399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11716__A (.DIODE(_05399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11234__A (.DIODE(_05399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13549__A0 (.DIODE(_05400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13413__A0 (.DIODE(_05400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13345__A0 (.DIODE(_05400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13277__A0 (.DIODE(_05400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13004__A0 (.DIODE(_05400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12732__A0 (.DIODE(_05400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12359__A0 (.DIODE(_05400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12077__A0 (.DIODE(_05400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11802__A0 (.DIODE(_05400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11235__A0 (.DIODE(_05400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11241__B2 (.DIODE(_05405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11255__B1 (.DIODE(_05419_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14070__A1 (.DIODE(_05423_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12583__A (.DIODE(_05423_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11719__A (.DIODE(_05423_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11259__A (.DIODE(_05423_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13551__A0 (.DIODE(_05424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13415__A0 (.DIODE(_05424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13347__A0 (.DIODE(_05424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13279__A0 (.DIODE(_05424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13006__A0 (.DIODE(_05424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12734__A0 (.DIODE(_05424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12361__A0 (.DIODE(_05424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12079__A0 (.DIODE(_05424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11804__A0 (.DIODE(_05424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11260__A0 (.DIODE(_05424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11265__B2 (.DIODE(_05428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11284__D_N (.DIODE(_05447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14072__A1 (.DIODE(_05451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12586__A (.DIODE(_05451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11722__A (.DIODE(_05451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11288__A (.DIODE(_05451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13553__A0 (.DIODE(_05452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13417__A0 (.DIODE(_05452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13349__A0 (.DIODE(_05452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13281__A0 (.DIODE(_05452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13008__A0 (.DIODE(_05452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12736__A0 (.DIODE(_05452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12363__A0 (.DIODE(_05452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12081__A0 (.DIODE(_05452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11806__A0 (.DIODE(_05452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11289__A0 (.DIODE(_05452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11296__B2 (.DIODE(_05458_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11311__C1 (.DIODE(_05473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14074__A1 (.DIODE(_05476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12589__A (.DIODE(_05476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11725__A (.DIODE(_05476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11314__A (.DIODE(_05476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13555__A0 (.DIODE(_05477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13419__A0 (.DIODE(_05477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13351__A0 (.DIODE(_05477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13283__A0 (.DIODE(_05477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13010__A0 (.DIODE(_05477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12738__A0 (.DIODE(_05477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12365__A0 (.DIODE(_05477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12083__A0 (.DIODE(_05477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11808__A0 (.DIODE(_05477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11315__A0 (.DIODE(_05477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11350__A2 (.DIODE(_05483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11329__B2 (.DIODE(_05485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11350__A4 (.DIODE(_05509_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14077__A1 (.DIODE(_05513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12592__A (.DIODE(_05513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11728__A (.DIODE(_05513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11352__A (.DIODE(_05513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13558__A0 (.DIODE(_05514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13422__A0 (.DIODE(_05514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13354__A0 (.DIODE(_05514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13286__A0 (.DIODE(_05514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13013__A0 (.DIODE(_05514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12741__A0 (.DIODE(_05514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12368__A0 (.DIODE(_05514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12086__A0 (.DIODE(_05514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11811__A0 (.DIODE(_05514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11354__A0 (.DIODE(_05514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11611__S (.DIODE(_05515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11582__S (.DIODE(_05515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11554__S (.DIODE(_05515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11529__S (.DIODE(_05515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11504__S (.DIODE(_05515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11479__S (.DIODE(_05515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11442__S (.DIODE(_05515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11411__S (.DIODE(_05515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11381__S (.DIODE(_05515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11354__S (.DIODE(_05515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11365__B2 (.DIODE(_05525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11377__D1 (.DIODE(_05537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13560__A0 (.DIODE(_05541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13424__A0 (.DIODE(_05541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13356__A0 (.DIODE(_05541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13288__A0 (.DIODE(_05541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13015__A0 (.DIODE(_05541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12743__A0 (.DIODE(_05541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12370__A0 (.DIODE(_05541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12088__A0 (.DIODE(_05541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11813__A0 (.DIODE(_05541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11381__A0 (.DIODE(_05541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11406__C1 (.DIODE(_05565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13562__A0 (.DIODE(_05570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13426__A0 (.DIODE(_05570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13358__A0 (.DIODE(_05570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13290__A0 (.DIODE(_05570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13017__A0 (.DIODE(_05570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12745__A0 (.DIODE(_05570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12372__A0 (.DIODE(_05570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12090__A0 (.DIODE(_05570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11815__A0 (.DIODE(_05570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11411__A0 (.DIODE(_05570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11437__B1 (.DIODE(_05591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11436__A2 (.DIODE(_05593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14083__A1 (.DIODE(_05599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12602__A (.DIODE(_05599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11738__A (.DIODE(_05599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11441__A (.DIODE(_05599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13564__A0 (.DIODE(_05600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13428__A0 (.DIODE(_05600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13360__A0 (.DIODE(_05600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13292__A0 (.DIODE(_05600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13019__A0 (.DIODE(_05600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12747__A0 (.DIODE(_05600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12374__A0 (.DIODE(_05600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12092__A0 (.DIODE(_05600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11817__A0 (.DIODE(_05600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11442__A0 (.DIODE(_05600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11573__A2 (.DIODE(_05613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11457__B (.DIODE(_05613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11456__B (.DIODE(_05613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11474__A3 (.DIODE(_05619_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11471__B2 (.DIODE(_05628_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13566__A0 (.DIODE(_05636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13430__A0 (.DIODE(_05636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13362__A0 (.DIODE(_05636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13294__A0 (.DIODE(_05636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13021__A0 (.DIODE(_05636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12749__A0 (.DIODE(_05636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12376__A0 (.DIODE(_05636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12094__A0 (.DIODE(_05636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11819__A0 (.DIODE(_05636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11479__A0 (.DIODE(_05636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11499__C1 (.DIODE(_05655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14087__A1 (.DIODE(_05659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12608__A (.DIODE(_05659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11744__A (.DIODE(_05659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11503__A (.DIODE(_05659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13568__A0 (.DIODE(_05660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13432__A0 (.DIODE(_05660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13364__A0 (.DIODE(_05660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13296__A0 (.DIODE(_05660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13023__A0 (.DIODE(_05660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12751__A0 (.DIODE(_05660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12378__A0 (.DIODE(_05660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12096__A0 (.DIODE(_05660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11821__A0 (.DIODE(_05660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11504__A0 (.DIODE(_05660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11524__A1 (.DIODE(_05668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11524__A2 (.DIODE(_05673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13570__A0 (.DIODE(_05684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13434__A0 (.DIODE(_05684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13366__A0 (.DIODE(_05684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13298__A0 (.DIODE(_05684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13025__A0 (.DIODE(_05684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12753__A0 (.DIODE(_05684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12380__A0 (.DIODE(_05684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12098__A0 (.DIODE(_05684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11823__A0 (.DIODE(_05684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11529__A0 (.DIODE(_05684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11552__A1 (.DIODE(_05697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14091__A1 (.DIODE(_05707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12614__A (.DIODE(_05707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11750__A (.DIODE(_05707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11553__A (.DIODE(_05707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13572__A0 (.DIODE(_05708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13436__A0 (.DIODE(_05708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13368__A0 (.DIODE(_05708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13300__A0 (.DIODE(_05708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13027__A0 (.DIODE(_05708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12755__A0 (.DIODE(_05708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12382__A0 (.DIODE(_05708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12100__A0 (.DIODE(_05708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11825__A0 (.DIODE(_05708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11554__A0 (.DIODE(_05708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11577__C1 (.DIODE(_05730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14093__A1 (.DIODE(_05734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12617__A (.DIODE(_05734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11753__A (.DIODE(_05734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11581__A (.DIODE(_05734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13574__A0 (.DIODE(_05735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13438__A0 (.DIODE(_05735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13370__A0 (.DIODE(_05735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13302__A0 (.DIODE(_05735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13029__A0 (.DIODE(_05735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12757__A0 (.DIODE(_05735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12384__A0 (.DIODE(_05735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12102__A0 (.DIODE(_05735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11827__A0 (.DIODE(_05735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11582__A0 (.DIODE(_05735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11609__A1 (.DIODE(_05751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13576__A0 (.DIODE(_05763_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13440__A0 (.DIODE(_05763_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13372__A0 (.DIODE(_05763_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13304__A0 (.DIODE(_05763_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13031__A0 (.DIODE(_05763_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12759__A0 (.DIODE(_05763_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12386__A0 (.DIODE(_05763_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12104__A0 (.DIODE(_05763_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11829__A0 (.DIODE(_05763_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11611__A0 (.DIODE(_05763_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11630__B2 (.DIODE(_05779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13578__A0 (.DIODE(_05787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13442__A0 (.DIODE(_05787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13374__A0 (.DIODE(_05787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13306__A0 (.DIODE(_05787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13033__A0 (.DIODE(_05787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12761__A0 (.DIODE(_05787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12388__A0 (.DIODE(_05787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12106__A0 (.DIODE(_05787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11831__A0 (.DIODE(_05787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11636__A0 (.DIODE(_05787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11652__B2 (.DIODE(_05802_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14099__A1 (.DIODE(_05810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12626__A (.DIODE(_05810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11762__A (.DIODE(_05810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11660__A (.DIODE(_05810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13580__A0 (.DIODE(_05811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13444__A0 (.DIODE(_05811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13376__A0 (.DIODE(_05811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13308__A0 (.DIODE(_05811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13035__A0 (.DIODE(_05811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12763__A0 (.DIODE(_05811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12390__A0 (.DIODE(_05811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12108__A0 (.DIODE(_05811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11833__A0 (.DIODE(_05811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11661__A0 (.DIODE(_05811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13652__A0 (.DIODE(_05813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12463__A1 (.DIODE(_05813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12395__A1 (.DIODE(_05813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12258__A1 (.DIODE(_05813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12189__A1 (.DIODE(_05813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12121__A1 (.DIODE(_05813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11975__A1 (.DIODE(_05813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11907__A1 (.DIODE(_05813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11838__A1 (.DIODE(_05813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11668__A1 (.DIODE(_05813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11763__S (.DIODE(_05816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11760__S (.DIODE(_05816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11729__A (.DIODE(_05816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11698__A (.DIODE(_05816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11667__A (.DIODE(_05816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11695__S (.DIODE(_05817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11692__S (.DIODE(_05817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11689__S (.DIODE(_05817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11686__S (.DIODE(_05817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11683__S (.DIODE(_05817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11680__S (.DIODE(_05817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11677__S (.DIODE(_05817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11674__S (.DIODE(_05817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11671__S (.DIODE(_05817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11668__S (.DIODE(_05817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13654__A0 (.DIODE(_05819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12465__A1 (.DIODE(_05819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12397__A1 (.DIODE(_05819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12260__A1 (.DIODE(_05819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12191__A1 (.DIODE(_05819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12123__A1 (.DIODE(_05819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11977__A1 (.DIODE(_05819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11909__A1 (.DIODE(_05819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11840__A1 (.DIODE(_05819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11671__A1 (.DIODE(_05819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13656__A0 (.DIODE(_05821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12467__A1 (.DIODE(_05821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12399__A1 (.DIODE(_05821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12262__A1 (.DIODE(_05821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12193__A1 (.DIODE(_05821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12125__A1 (.DIODE(_05821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11979__A1 (.DIODE(_05821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11911__A1 (.DIODE(_05821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11842__A1 (.DIODE(_05821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11674__A1 (.DIODE(_05821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13658__A0 (.DIODE(_05823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12469__A1 (.DIODE(_05823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12401__A1 (.DIODE(_05823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12264__A1 (.DIODE(_05823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12195__A1 (.DIODE(_05823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12127__A1 (.DIODE(_05823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11981__A1 (.DIODE(_05823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11913__A1 (.DIODE(_05823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11844__A1 (.DIODE(_05823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11677__A1 (.DIODE(_05823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13660__A0 (.DIODE(_05825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12471__A1 (.DIODE(_05825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12403__A1 (.DIODE(_05825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12266__A1 (.DIODE(_05825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12197__A1 (.DIODE(_05825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12129__A1 (.DIODE(_05825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11983__A1 (.DIODE(_05825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11915__A1 (.DIODE(_05825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11846__A1 (.DIODE(_05825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11680__A1 (.DIODE(_05825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13662__A0 (.DIODE(_05827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12473__A1 (.DIODE(_05827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12405__A1 (.DIODE(_05827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12268__A1 (.DIODE(_05827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12199__A1 (.DIODE(_05827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12131__A1 (.DIODE(_05827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11985__A1 (.DIODE(_05827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11917__A1 (.DIODE(_05827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11848__A1 (.DIODE(_05827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11683__A1 (.DIODE(_05827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13664__A0 (.DIODE(_05829_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12475__A1 (.DIODE(_05829_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12407__A1 (.DIODE(_05829_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12270__A1 (.DIODE(_05829_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12201__A1 (.DIODE(_05829_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12133__A1 (.DIODE(_05829_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11987__A1 (.DIODE(_05829_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11919__A1 (.DIODE(_05829_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11850__A1 (.DIODE(_05829_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11686__A1 (.DIODE(_05829_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13666__A0 (.DIODE(_05831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12477__A1 (.DIODE(_05831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12409__A1 (.DIODE(_05831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12272__A1 (.DIODE(_05831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12203__A1 (.DIODE(_05831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12135__A1 (.DIODE(_05831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11989__A1 (.DIODE(_05831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11921__A1 (.DIODE(_05831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11852__A1 (.DIODE(_05831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11689__A1 (.DIODE(_05831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13668__A0 (.DIODE(_05833_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12479__A1 (.DIODE(_05833_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12411__A1 (.DIODE(_05833_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12274__A1 (.DIODE(_05833_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12205__A1 (.DIODE(_05833_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12137__A1 (.DIODE(_05833_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11991__A1 (.DIODE(_05833_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11923__A1 (.DIODE(_05833_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11854__A1 (.DIODE(_05833_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11692__A1 (.DIODE(_05833_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13670__A0 (.DIODE(_05835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12481__A1 (.DIODE(_05835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12413__A1 (.DIODE(_05835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12276__A1 (.DIODE(_05835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12207__A1 (.DIODE(_05835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12139__A1 (.DIODE(_05835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11993__A1 (.DIODE(_05835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11925__A1 (.DIODE(_05835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11856__A1 (.DIODE(_05835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11695__A1 (.DIODE(_05835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13673__A0 (.DIODE(_05837_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12484__A1 (.DIODE(_05837_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12416__A1 (.DIODE(_05837_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12279__A1 (.DIODE(_05837_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12210__A1 (.DIODE(_05837_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12142__A1 (.DIODE(_05837_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11996__A1 (.DIODE(_05837_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11928__A1 (.DIODE(_05837_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11859__A1 (.DIODE(_05837_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11699__A1 (.DIODE(_05837_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11726__S (.DIODE(_05838_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11723__S (.DIODE(_05838_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11720__S (.DIODE(_05838_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11717__S (.DIODE(_05838_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11714__S (.DIODE(_05838_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11711__S (.DIODE(_05838_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11708__S (.DIODE(_05838_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11705__S (.DIODE(_05838_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11702__S (.DIODE(_05838_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11699__S (.DIODE(_05838_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13675__A0 (.DIODE(_05840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12486__A1 (.DIODE(_05840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12418__A1 (.DIODE(_05840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12281__A1 (.DIODE(_05840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12212__A1 (.DIODE(_05840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12144__A1 (.DIODE(_05840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11998__A1 (.DIODE(_05840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11930__A1 (.DIODE(_05840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11861__A1 (.DIODE(_05840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11702__A1 (.DIODE(_05840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13677__A0 (.DIODE(_05842_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12488__A1 (.DIODE(_05842_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12420__A1 (.DIODE(_05842_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12283__A1 (.DIODE(_05842_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12214__A1 (.DIODE(_05842_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12146__A1 (.DIODE(_05842_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12000__A1 (.DIODE(_05842_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11932__A1 (.DIODE(_05842_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11863__A1 (.DIODE(_05842_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11705__A1 (.DIODE(_05842_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13679__A0 (.DIODE(_05844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12490__A1 (.DIODE(_05844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12422__A1 (.DIODE(_05844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12285__A1 (.DIODE(_05844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12216__A1 (.DIODE(_05844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12148__A1 (.DIODE(_05844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12002__A1 (.DIODE(_05844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11934__A1 (.DIODE(_05844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11865__A1 (.DIODE(_05844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11708__A1 (.DIODE(_05844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13681__A0 (.DIODE(_05846_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12492__A1 (.DIODE(_05846_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12424__A1 (.DIODE(_05846_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12287__A1 (.DIODE(_05846_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12218__A1 (.DIODE(_05846_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12150__A1 (.DIODE(_05846_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12004__A1 (.DIODE(_05846_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11936__A1 (.DIODE(_05846_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11867__A1 (.DIODE(_05846_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11711__A1 (.DIODE(_05846_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13683__A0 (.DIODE(_05848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12494__A1 (.DIODE(_05848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12426__A1 (.DIODE(_05848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12289__A1 (.DIODE(_05848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12220__A1 (.DIODE(_05848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12152__A1 (.DIODE(_05848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12006__A1 (.DIODE(_05848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11938__A1 (.DIODE(_05848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11869__A1 (.DIODE(_05848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11714__A1 (.DIODE(_05848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13685__A0 (.DIODE(_05850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12496__A1 (.DIODE(_05850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12428__A1 (.DIODE(_05850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12291__A1 (.DIODE(_05850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12222__A1 (.DIODE(_05850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12154__A1 (.DIODE(_05850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12008__A1 (.DIODE(_05850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11940__A1 (.DIODE(_05850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11871__A1 (.DIODE(_05850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11717__A1 (.DIODE(_05850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13687__A0 (.DIODE(_05852_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12498__A1 (.DIODE(_05852_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12430__A1 (.DIODE(_05852_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12293__A1 (.DIODE(_05852_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12224__A1 (.DIODE(_05852_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12156__A1 (.DIODE(_05852_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12010__A1 (.DIODE(_05852_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11942__A1 (.DIODE(_05852_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11873__A1 (.DIODE(_05852_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11720__A1 (.DIODE(_05852_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13689__A0 (.DIODE(_05854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12500__A1 (.DIODE(_05854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12432__A1 (.DIODE(_05854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12295__A1 (.DIODE(_05854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12226__A1 (.DIODE(_05854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12158__A1 (.DIODE(_05854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12012__A1 (.DIODE(_05854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11944__A1 (.DIODE(_05854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11875__A1 (.DIODE(_05854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11723__A1 (.DIODE(_05854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13691__A0 (.DIODE(_05856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12502__A1 (.DIODE(_05856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12434__A1 (.DIODE(_05856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12297__A1 (.DIODE(_05856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12228__A1 (.DIODE(_05856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12160__A1 (.DIODE(_05856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12014__A1 (.DIODE(_05856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11946__A1 (.DIODE(_05856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11877__A1 (.DIODE(_05856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11726__A1 (.DIODE(_05856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13694__A0 (.DIODE(_05858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12505__A1 (.DIODE(_05858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12437__A1 (.DIODE(_05858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12300__A1 (.DIODE(_05858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12231__A1 (.DIODE(_05858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12163__A1 (.DIODE(_05858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12017__A1 (.DIODE(_05858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11949__A1 (.DIODE(_05858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11880__A1 (.DIODE(_05858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11730__A1 (.DIODE(_05858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11757__S (.DIODE(_05859_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11754__S (.DIODE(_05859_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11751__S (.DIODE(_05859_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11748__S (.DIODE(_05859_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11745__S (.DIODE(_05859_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11742__S (.DIODE(_05859_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11739__S (.DIODE(_05859_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11736__S (.DIODE(_05859_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11733__S (.DIODE(_05859_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11730__S (.DIODE(_05859_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13696__A0 (.DIODE(_05861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12507__A1 (.DIODE(_05861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12439__A1 (.DIODE(_05861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12302__A1 (.DIODE(_05861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12233__A1 (.DIODE(_05861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12165__A1 (.DIODE(_05861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12019__A1 (.DIODE(_05861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11951__A1 (.DIODE(_05861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11882__A1 (.DIODE(_05861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11733__A1 (.DIODE(_05861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13698__A0 (.DIODE(_05863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12509__A1 (.DIODE(_05863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12441__A1 (.DIODE(_05863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12304__A1 (.DIODE(_05863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12235__A1 (.DIODE(_05863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12167__A1 (.DIODE(_05863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12021__A1 (.DIODE(_05863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11953__A1 (.DIODE(_05863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11884__A1 (.DIODE(_05863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11736__A1 (.DIODE(_05863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13700__A0 (.DIODE(_05865_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12511__A1 (.DIODE(_05865_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12443__A1 (.DIODE(_05865_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12306__A1 (.DIODE(_05865_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12237__A1 (.DIODE(_05865_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12169__A1 (.DIODE(_05865_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12023__A1 (.DIODE(_05865_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11955__A1 (.DIODE(_05865_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11886__A1 (.DIODE(_05865_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11739__A1 (.DIODE(_05865_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13702__A0 (.DIODE(_05867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12513__A1 (.DIODE(_05867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12445__A1 (.DIODE(_05867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12308__A1 (.DIODE(_05867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12239__A1 (.DIODE(_05867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12171__A1 (.DIODE(_05867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12025__A1 (.DIODE(_05867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11957__A1 (.DIODE(_05867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11888__A1 (.DIODE(_05867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11742__A1 (.DIODE(_05867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13704__A0 (.DIODE(_05869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12515__A1 (.DIODE(_05869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12447__A1 (.DIODE(_05869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12310__A1 (.DIODE(_05869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12241__A1 (.DIODE(_05869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12173__A1 (.DIODE(_05869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12027__A1 (.DIODE(_05869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11959__A1 (.DIODE(_05869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11890__A1 (.DIODE(_05869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11745__A1 (.DIODE(_05869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13706__A0 (.DIODE(_05871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12517__A1 (.DIODE(_05871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12449__A1 (.DIODE(_05871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12312__A1 (.DIODE(_05871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12243__A1 (.DIODE(_05871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12175__A1 (.DIODE(_05871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12029__A1 (.DIODE(_05871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11961__A1 (.DIODE(_05871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11892__A1 (.DIODE(_05871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11748__A1 (.DIODE(_05871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13708__A0 (.DIODE(_05873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12519__A1 (.DIODE(_05873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12451__A1 (.DIODE(_05873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12314__A1 (.DIODE(_05873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12245__A1 (.DIODE(_05873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12177__A1 (.DIODE(_05873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12031__A1 (.DIODE(_05873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11963__A1 (.DIODE(_05873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11894__A1 (.DIODE(_05873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11751__A1 (.DIODE(_05873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13710__A0 (.DIODE(_05875_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12521__A1 (.DIODE(_05875_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12453__A1 (.DIODE(_05875_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12316__A1 (.DIODE(_05875_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12247__A1 (.DIODE(_05875_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12179__A1 (.DIODE(_05875_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12033__A1 (.DIODE(_05875_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11965__A1 (.DIODE(_05875_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11896__A1 (.DIODE(_05875_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11754__A1 (.DIODE(_05875_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13712__A0 (.DIODE(_05877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12523__A1 (.DIODE(_05877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12455__A1 (.DIODE(_05877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12318__A1 (.DIODE(_05877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12249__A1 (.DIODE(_05877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12181__A1 (.DIODE(_05877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12035__A1 (.DIODE(_05877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11967__A1 (.DIODE(_05877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11898__A1 (.DIODE(_05877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11757__A1 (.DIODE(_05877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13714__A0 (.DIODE(_05879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12525__A1 (.DIODE(_05879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12457__A1 (.DIODE(_05879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12320__A1 (.DIODE(_05879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12251__A1 (.DIODE(_05879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12183__A1 (.DIODE(_05879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12037__A1 (.DIODE(_05879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11969__A1 (.DIODE(_05879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11900__A1 (.DIODE(_05879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11760__A1 (.DIODE(_05879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11833__S (.DIODE(_05885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11831__S (.DIODE(_05885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11810__A (.DIODE(_05885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11789__A (.DIODE(_05885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11768__A (.DIODE(_05885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11787__S (.DIODE(_05886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11785__S (.DIODE(_05886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11783__S (.DIODE(_05886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11781__S (.DIODE(_05886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11779__S (.DIODE(_05886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11777__S (.DIODE(_05886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11775__S (.DIODE(_05886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11773__S (.DIODE(_05886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11771__S (.DIODE(_05886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11769__S (.DIODE(_05886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11808__S (.DIODE(_05897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11806__S (.DIODE(_05897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11804__S (.DIODE(_05897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11802__S (.DIODE(_05897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11800__S (.DIODE(_05897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11798__S (.DIODE(_05897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11796__S (.DIODE(_05897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11794__S (.DIODE(_05897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11792__S (.DIODE(_05897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11790__S (.DIODE(_05897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11829__S (.DIODE(_05908_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11827__S (.DIODE(_05908_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11825__S (.DIODE(_05908_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11823__S (.DIODE(_05908_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11821__S (.DIODE(_05908_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11819__S (.DIODE(_05908_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11817__S (.DIODE(_05908_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11815__S (.DIODE(_05908_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11813__S (.DIODE(_05908_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11811__S (.DIODE(_05908_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11902__S (.DIODE(_05922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11900__S (.DIODE(_05922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11879__A (.DIODE(_05922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11858__A (.DIODE(_05922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11837__A (.DIODE(_05922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11856__S (.DIODE(_05923_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11854__S (.DIODE(_05923_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11852__S (.DIODE(_05923_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11850__S (.DIODE(_05923_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11848__S (.DIODE(_05923_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11846__S (.DIODE(_05923_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11844__S (.DIODE(_05923_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11842__S (.DIODE(_05923_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11840__S (.DIODE(_05923_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11838__S (.DIODE(_05923_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11877__S (.DIODE(_05934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11875__S (.DIODE(_05934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11873__S (.DIODE(_05934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11871__S (.DIODE(_05934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11869__S (.DIODE(_05934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11867__S (.DIODE(_05934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11865__S (.DIODE(_05934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11863__S (.DIODE(_05934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11861__S (.DIODE(_05934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11859__S (.DIODE(_05934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11898__S (.DIODE(_05945_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11896__S (.DIODE(_05945_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11894__S (.DIODE(_05945_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11892__S (.DIODE(_05945_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11890__S (.DIODE(_05945_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11888__S (.DIODE(_05945_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11886__S (.DIODE(_05945_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11884__S (.DIODE(_05945_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11882__S (.DIODE(_05945_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11880__S (.DIODE(_05945_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11971__S (.DIODE(_05959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11969__S (.DIODE(_05959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11948__A (.DIODE(_05959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11927__A (.DIODE(_05959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11906__A (.DIODE(_05959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11925__S (.DIODE(_05960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11923__S (.DIODE(_05960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11921__S (.DIODE(_05960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11919__S (.DIODE(_05960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11917__S (.DIODE(_05960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11915__S (.DIODE(_05960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11913__S (.DIODE(_05960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11911__S (.DIODE(_05960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11909__S (.DIODE(_05960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11907__S (.DIODE(_05960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11946__S (.DIODE(_05971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11944__S (.DIODE(_05971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11942__S (.DIODE(_05971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11940__S (.DIODE(_05971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11938__S (.DIODE(_05971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11936__S (.DIODE(_05971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11934__S (.DIODE(_05971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11932__S (.DIODE(_05971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11930__S (.DIODE(_05971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11928__S (.DIODE(_05971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11967__S (.DIODE(_05982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11965__S (.DIODE(_05982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11963__S (.DIODE(_05982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11961__S (.DIODE(_05982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11959__S (.DIODE(_05982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11957__S (.DIODE(_05982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11955__S (.DIODE(_05982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11953__S (.DIODE(_05982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11951__S (.DIODE(_05982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11949__S (.DIODE(_05982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12039__S (.DIODE(_05995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12037__S (.DIODE(_05995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12016__A (.DIODE(_05995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11995__A (.DIODE(_05995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11974__A (.DIODE(_05995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11993__S (.DIODE(_05996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11991__S (.DIODE(_05996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11989__S (.DIODE(_05996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11987__S (.DIODE(_05996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11985__S (.DIODE(_05996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11983__S (.DIODE(_05996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11981__S (.DIODE(_05996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11979__S (.DIODE(_05996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11977__S (.DIODE(_05996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11975__S (.DIODE(_05996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12014__S (.DIODE(_06007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12012__S (.DIODE(_06007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12010__S (.DIODE(_06007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12008__S (.DIODE(_06007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12006__S (.DIODE(_06007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12004__S (.DIODE(_06007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12002__S (.DIODE(_06007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12000__S (.DIODE(_06007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11998__S (.DIODE(_06007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11996__S (.DIODE(_06007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12035__S (.DIODE(_06018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12033__S (.DIODE(_06018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12031__S (.DIODE(_06018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12029__S (.DIODE(_06018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12027__S (.DIODE(_06018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12025__S (.DIODE(_06018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12023__S (.DIODE(_06018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12021__S (.DIODE(_06018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12019__S (.DIODE(_06018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12017__S (.DIODE(_06018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12108__S (.DIODE(_06032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12106__S (.DIODE(_06032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12085__A (.DIODE(_06032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12064__A (.DIODE(_06032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12043__A (.DIODE(_06032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12062__S (.DIODE(_06033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12060__S (.DIODE(_06033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12058__S (.DIODE(_06033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12056__S (.DIODE(_06033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12054__S (.DIODE(_06033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12052__S (.DIODE(_06033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12050__S (.DIODE(_06033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12048__S (.DIODE(_06033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12046__S (.DIODE(_06033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12044__S (.DIODE(_06033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12083__S (.DIODE(_06044_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12081__S (.DIODE(_06044_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12079__S (.DIODE(_06044_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12077__S (.DIODE(_06044_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12075__S (.DIODE(_06044_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12073__S (.DIODE(_06044_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12071__S (.DIODE(_06044_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12069__S (.DIODE(_06044_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12067__S (.DIODE(_06044_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12065__S (.DIODE(_06044_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12104__S (.DIODE(_06055_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12102__S (.DIODE(_06055_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12100__S (.DIODE(_06055_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12098__S (.DIODE(_06055_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12096__S (.DIODE(_06055_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12094__S (.DIODE(_06055_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12092__S (.DIODE(_06055_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12090__S (.DIODE(_06055_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12088__S (.DIODE(_06055_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12086__S (.DIODE(_06055_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12830__A (.DIODE(_06068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12828__A (.DIODE(_06068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12826__A (.DIODE(_06068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12805__A (.DIODE(_06068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12784__A (.DIODE(_06068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12111__A (.DIODE(_06068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13880__A (.DIODE(_06069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13869__A (.DIODE(_06069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13858__A (.DIODE(_06069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13847__A (.DIODE(_06069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13836__A (.DIODE(_06069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13825__A (.DIODE(_06069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13814__A (.DIODE(_06069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13803__A (.DIODE(_06069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13792__A (.DIODE(_06069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12113__A (.DIODE(_06069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13791__A (.DIODE(_06070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13790__A (.DIODE(_06070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13789__A (.DIODE(_06070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13788__A (.DIODE(_06070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13787__A (.DIODE(_06070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13786__A (.DIODE(_06070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12765__A (.DIODE(_06070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12116__A (.DIODE(_06070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12115__A (.DIODE(_06070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12114__A (.DIODE(_06070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12185__S (.DIODE(_06073_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12183__S (.DIODE(_06073_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12162__A (.DIODE(_06073_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12141__A (.DIODE(_06073_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12120__A (.DIODE(_06073_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12139__S (.DIODE(_06074_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12137__S (.DIODE(_06074_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12135__S (.DIODE(_06074_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12133__S (.DIODE(_06074_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12131__S (.DIODE(_06074_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12129__S (.DIODE(_06074_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12127__S (.DIODE(_06074_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12125__S (.DIODE(_06074_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12123__S (.DIODE(_06074_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12121__S (.DIODE(_06074_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12160__S (.DIODE(_06085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12158__S (.DIODE(_06085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12156__S (.DIODE(_06085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12154__S (.DIODE(_06085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12152__S (.DIODE(_06085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12150__S (.DIODE(_06085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12148__S (.DIODE(_06085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12146__S (.DIODE(_06085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12144__S (.DIODE(_06085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12142__S (.DIODE(_06085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12181__S (.DIODE(_06096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12179__S (.DIODE(_06096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12177__S (.DIODE(_06096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12175__S (.DIODE(_06096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12173__S (.DIODE(_06096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12171__S (.DIODE(_06096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12169__S (.DIODE(_06096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12167__S (.DIODE(_06096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12165__S (.DIODE(_06096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12163__S (.DIODE(_06096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12253__S (.DIODE(_06109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12251__S (.DIODE(_06109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12230__A (.DIODE(_06109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12209__A (.DIODE(_06109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12188__A (.DIODE(_06109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12207__S (.DIODE(_06110_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12205__S (.DIODE(_06110_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12203__S (.DIODE(_06110_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12201__S (.DIODE(_06110_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12199__S (.DIODE(_06110_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12197__S (.DIODE(_06110_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12195__S (.DIODE(_06110_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12193__S (.DIODE(_06110_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12191__S (.DIODE(_06110_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12189__S (.DIODE(_06110_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12228__S (.DIODE(_06121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12226__S (.DIODE(_06121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12224__S (.DIODE(_06121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12222__S (.DIODE(_06121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12220__S (.DIODE(_06121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12218__S (.DIODE(_06121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12216__S (.DIODE(_06121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12214__S (.DIODE(_06121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12212__S (.DIODE(_06121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12210__S (.DIODE(_06121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12249__S (.DIODE(_06132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12247__S (.DIODE(_06132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12245__S (.DIODE(_06132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12243__S (.DIODE(_06132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12241__S (.DIODE(_06132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12239__S (.DIODE(_06132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12237__S (.DIODE(_06132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12235__S (.DIODE(_06132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12233__S (.DIODE(_06132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12231__S (.DIODE(_06132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12276__S (.DIODE(_06147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12274__S (.DIODE(_06147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12272__S (.DIODE(_06147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12270__S (.DIODE(_06147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12268__S (.DIODE(_06147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12266__S (.DIODE(_06147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12264__S (.DIODE(_06147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12262__S (.DIODE(_06147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12260__S (.DIODE(_06147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12258__S (.DIODE(_06147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12297__S (.DIODE(_06158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12295__S (.DIODE(_06158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12293__S (.DIODE(_06158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12291__S (.DIODE(_06158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12289__S (.DIODE(_06158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12287__S (.DIODE(_06158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12285__S (.DIODE(_06158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12283__S (.DIODE(_06158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12281__S (.DIODE(_06158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12279__S (.DIODE(_06158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12318__S (.DIODE(_06169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12316__S (.DIODE(_06169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12314__S (.DIODE(_06169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12312__S (.DIODE(_06169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12310__S (.DIODE(_06169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12308__S (.DIODE(_06169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12306__S (.DIODE(_06169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12304__S (.DIODE(_06169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12302__S (.DIODE(_06169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12300__S (.DIODE(_06169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12390__S (.DIODE(_06182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12388__S (.DIODE(_06182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12367__A (.DIODE(_06182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12346__A (.DIODE(_06182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12325__A (.DIODE(_06182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12344__S (.DIODE(_06183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12342__S (.DIODE(_06183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12340__S (.DIODE(_06183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12338__S (.DIODE(_06183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12336__S (.DIODE(_06183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12334__S (.DIODE(_06183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12332__S (.DIODE(_06183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12330__S (.DIODE(_06183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12328__S (.DIODE(_06183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12326__S (.DIODE(_06183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12365__S (.DIODE(_06194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12363__S (.DIODE(_06194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12361__S (.DIODE(_06194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12359__S (.DIODE(_06194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12357__S (.DIODE(_06194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12355__S (.DIODE(_06194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12353__S (.DIODE(_06194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12351__S (.DIODE(_06194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12349__S (.DIODE(_06194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12347__S (.DIODE(_06194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12386__S (.DIODE(_06205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12384__S (.DIODE(_06205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12382__S (.DIODE(_06205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12380__S (.DIODE(_06205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12378__S (.DIODE(_06205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12376__S (.DIODE(_06205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12374__S (.DIODE(_06205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12372__S (.DIODE(_06205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12370__S (.DIODE(_06205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12368__S (.DIODE(_06205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12413__S (.DIODE(_06220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12411__S (.DIODE(_06220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12409__S (.DIODE(_06220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12407__S (.DIODE(_06220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12405__S (.DIODE(_06220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12403__S (.DIODE(_06220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12401__S (.DIODE(_06220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12399__S (.DIODE(_06220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12397__S (.DIODE(_06220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12395__S (.DIODE(_06220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12434__S (.DIODE(_06231_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12432__S (.DIODE(_06231_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12430__S (.DIODE(_06231_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12428__S (.DIODE(_06231_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12426__S (.DIODE(_06231_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12424__S (.DIODE(_06231_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12422__S (.DIODE(_06231_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12420__S (.DIODE(_06231_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12418__S (.DIODE(_06231_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12416__S (.DIODE(_06231_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12455__S (.DIODE(_06242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12453__S (.DIODE(_06242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12451__S (.DIODE(_06242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12449__S (.DIODE(_06242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12447__S (.DIODE(_06242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12445__S (.DIODE(_06242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12443__S (.DIODE(_06242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12441__S (.DIODE(_06242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12439__S (.DIODE(_06242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12437__S (.DIODE(_06242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12481__S (.DIODE(_06256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12479__S (.DIODE(_06256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12477__S (.DIODE(_06256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12475__S (.DIODE(_06256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12473__S (.DIODE(_06256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12471__S (.DIODE(_06256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12469__S (.DIODE(_06256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12467__S (.DIODE(_06256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12465__S (.DIODE(_06256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12463__S (.DIODE(_06256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12502__S (.DIODE(_06267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12500__S (.DIODE(_06267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12498__S (.DIODE(_06267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12496__S (.DIODE(_06267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12494__S (.DIODE(_06267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12492__S (.DIODE(_06267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12490__S (.DIODE(_06267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12488__S (.DIODE(_06267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12486__S (.DIODE(_06267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12484__S (.DIODE(_06267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12523__S (.DIODE(_06278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12521__S (.DIODE(_06278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12519__S (.DIODE(_06278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12517__S (.DIODE(_06278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12515__S (.DIODE(_06278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12513__S (.DIODE(_06278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12511__S (.DIODE(_06278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12509__S (.DIODE(_06278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12507__S (.DIODE(_06278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12505__S (.DIODE(_06278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13720__A1 (.DIODE(_06291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13584__A1 (.DIODE(_06291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13448__A1 (.DIODE(_06291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13175__A1 (.DIODE(_06291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13107__A1 (.DIODE(_06291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13039__A1 (.DIODE(_06291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12902__A1 (.DIODE(_06291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12834__A1 (.DIODE(_06291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12631__A1 (.DIODE(_06291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12532__A1 (.DIODE(_06291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12627__S (.DIODE(_06292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12624__S (.DIODE(_06292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12593__A (.DIODE(_06292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12562__A (.DIODE(_06292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12531__A (.DIODE(_06292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12559__S (.DIODE(_06293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12556__S (.DIODE(_06293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12553__S (.DIODE(_06293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12550__S (.DIODE(_06293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12547__S (.DIODE(_06293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12544__S (.DIODE(_06293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12541__S (.DIODE(_06293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12538__S (.DIODE(_06293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12535__S (.DIODE(_06293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12532__S (.DIODE(_06293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13722__A1 (.DIODE(_06295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13586__A1 (.DIODE(_06295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13450__A1 (.DIODE(_06295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13177__A1 (.DIODE(_06295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13109__A1 (.DIODE(_06295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13041__A1 (.DIODE(_06295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12904__A1 (.DIODE(_06295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12836__A1 (.DIODE(_06295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12633__A1 (.DIODE(_06295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12535__A1 (.DIODE(_06295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13724__A1 (.DIODE(_06297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13588__A1 (.DIODE(_06297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13452__A1 (.DIODE(_06297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13179__A1 (.DIODE(_06297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13111__A1 (.DIODE(_06297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13043__A1 (.DIODE(_06297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12906__A1 (.DIODE(_06297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12838__A1 (.DIODE(_06297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12635__A1 (.DIODE(_06297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12538__A1 (.DIODE(_06297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13726__A1 (.DIODE(_06299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13590__A1 (.DIODE(_06299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13454__A1 (.DIODE(_06299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13181__A1 (.DIODE(_06299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13113__A1 (.DIODE(_06299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13045__A1 (.DIODE(_06299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12908__A1 (.DIODE(_06299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12840__A1 (.DIODE(_06299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12637__A1 (.DIODE(_06299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12541__A1 (.DIODE(_06299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13728__A1 (.DIODE(_06301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13592__A1 (.DIODE(_06301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13456__A1 (.DIODE(_06301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13183__A1 (.DIODE(_06301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13115__A1 (.DIODE(_06301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13047__A1 (.DIODE(_06301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12910__A1 (.DIODE(_06301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12842__A1 (.DIODE(_06301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12639__A1 (.DIODE(_06301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12544__A1 (.DIODE(_06301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13730__A1 (.DIODE(_06303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13594__A1 (.DIODE(_06303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13458__A1 (.DIODE(_06303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13185__A1 (.DIODE(_06303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13117__A1 (.DIODE(_06303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13049__A1 (.DIODE(_06303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12912__A1 (.DIODE(_06303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12844__A1 (.DIODE(_06303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12641__A1 (.DIODE(_06303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12547__A1 (.DIODE(_06303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13732__A1 (.DIODE(_06305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13596__A1 (.DIODE(_06305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13460__A1 (.DIODE(_06305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13187__A1 (.DIODE(_06305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13119__A1 (.DIODE(_06305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13051__A1 (.DIODE(_06305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12914__A1 (.DIODE(_06305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12846__A1 (.DIODE(_06305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12643__A1 (.DIODE(_06305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12550__A1 (.DIODE(_06305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13734__A1 (.DIODE(_06307_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13598__A1 (.DIODE(_06307_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13462__A1 (.DIODE(_06307_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13189__A1 (.DIODE(_06307_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13121__A1 (.DIODE(_06307_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13053__A1 (.DIODE(_06307_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12916__A1 (.DIODE(_06307_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12848__A1 (.DIODE(_06307_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12645__A1 (.DIODE(_06307_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12553__A1 (.DIODE(_06307_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13736__A1 (.DIODE(_06309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13600__A1 (.DIODE(_06309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13464__A1 (.DIODE(_06309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13191__A1 (.DIODE(_06309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13123__A1 (.DIODE(_06309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13055__A1 (.DIODE(_06309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12918__A1 (.DIODE(_06309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12850__A1 (.DIODE(_06309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12647__A1 (.DIODE(_06309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12556__A1 (.DIODE(_06309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13738__A1 (.DIODE(_06311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13602__A1 (.DIODE(_06311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13466__A1 (.DIODE(_06311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13193__A1 (.DIODE(_06311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13125__A1 (.DIODE(_06311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13057__A1 (.DIODE(_06311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12920__A1 (.DIODE(_06311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12852__A1 (.DIODE(_06311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12649__A1 (.DIODE(_06311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12559__A1 (.DIODE(_06311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13741__A1 (.DIODE(_06313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13605__A1 (.DIODE(_06313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13469__A1 (.DIODE(_06313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13196__A1 (.DIODE(_06313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13128__A1 (.DIODE(_06313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13060__A1 (.DIODE(_06313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12923__A1 (.DIODE(_06313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12855__A1 (.DIODE(_06313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12652__A1 (.DIODE(_06313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12563__A1 (.DIODE(_06313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12590__S (.DIODE(_06314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12587__S (.DIODE(_06314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12584__S (.DIODE(_06314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12581__S (.DIODE(_06314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12578__S (.DIODE(_06314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12575__S (.DIODE(_06314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12572__S (.DIODE(_06314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12569__S (.DIODE(_06314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12566__S (.DIODE(_06314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12563__S (.DIODE(_06314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13743__A1 (.DIODE(_06316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13607__A1 (.DIODE(_06316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13471__A1 (.DIODE(_06316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13198__A1 (.DIODE(_06316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13130__A1 (.DIODE(_06316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13062__A1 (.DIODE(_06316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12925__A1 (.DIODE(_06316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12857__A1 (.DIODE(_06316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12654__A1 (.DIODE(_06316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12566__A1 (.DIODE(_06316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13745__A1 (.DIODE(_06318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13609__A1 (.DIODE(_06318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13473__A1 (.DIODE(_06318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13200__A1 (.DIODE(_06318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13132__A1 (.DIODE(_06318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13064__A1 (.DIODE(_06318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12927__A1 (.DIODE(_06318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12859__A1 (.DIODE(_06318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12656__A1 (.DIODE(_06318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12569__A1 (.DIODE(_06318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13747__A1 (.DIODE(_06320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13611__A1 (.DIODE(_06320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13475__A1 (.DIODE(_06320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13202__A1 (.DIODE(_06320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13134__A1 (.DIODE(_06320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13066__A1 (.DIODE(_06320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12929__A1 (.DIODE(_06320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12861__A1 (.DIODE(_06320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12658__A1 (.DIODE(_06320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12572__A1 (.DIODE(_06320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13749__A1 (.DIODE(_06322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13613__A1 (.DIODE(_06322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13477__A1 (.DIODE(_06322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13204__A1 (.DIODE(_06322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13136__A1 (.DIODE(_06322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13068__A1 (.DIODE(_06322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12931__A1 (.DIODE(_06322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12863__A1 (.DIODE(_06322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12660__A1 (.DIODE(_06322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12575__A1 (.DIODE(_06322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13753__A1 (.DIODE(_06326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13617__A1 (.DIODE(_06326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13481__A1 (.DIODE(_06326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13208__A1 (.DIODE(_06326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13140__A1 (.DIODE(_06326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13072__A1 (.DIODE(_06326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12935__A1 (.DIODE(_06326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12867__A1 (.DIODE(_06326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12664__A1 (.DIODE(_06326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12581__A1 (.DIODE(_06326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13755__A1 (.DIODE(_06328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13619__A1 (.DIODE(_06328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13483__A1 (.DIODE(_06328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13210__A1 (.DIODE(_06328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13142__A1 (.DIODE(_06328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13074__A1 (.DIODE(_06328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12937__A1 (.DIODE(_06328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12869__A1 (.DIODE(_06328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12666__A1 (.DIODE(_06328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12584__A1 (.DIODE(_06328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13757__A1 (.DIODE(_06330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13621__A1 (.DIODE(_06330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13485__A1 (.DIODE(_06330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13212__A1 (.DIODE(_06330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13144__A1 (.DIODE(_06330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13076__A1 (.DIODE(_06330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12939__A1 (.DIODE(_06330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12871__A1 (.DIODE(_06330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12668__A1 (.DIODE(_06330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12587__A1 (.DIODE(_06330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13759__A1 (.DIODE(_06332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13623__A1 (.DIODE(_06332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13487__A1 (.DIODE(_06332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13214__A1 (.DIODE(_06332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13146__A1 (.DIODE(_06332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13078__A1 (.DIODE(_06332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12941__A1 (.DIODE(_06332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12873__A1 (.DIODE(_06332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12670__A1 (.DIODE(_06332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12590__A1 (.DIODE(_06332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13762__A1 (.DIODE(_06334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13626__A1 (.DIODE(_06334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13490__A1 (.DIODE(_06334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13217__A1 (.DIODE(_06334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13149__A1 (.DIODE(_06334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13081__A1 (.DIODE(_06334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12944__A1 (.DIODE(_06334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12876__A1 (.DIODE(_06334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12673__A1 (.DIODE(_06334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12594__A1 (.DIODE(_06334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12621__S (.DIODE(_06335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12618__S (.DIODE(_06335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12615__S (.DIODE(_06335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12612__S (.DIODE(_06335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12609__S (.DIODE(_06335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12606__S (.DIODE(_06335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12603__S (.DIODE(_06335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12600__S (.DIODE(_06335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12597__S (.DIODE(_06335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12594__S (.DIODE(_06335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13764__A1 (.DIODE(_06337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13628__A1 (.DIODE(_06337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13492__A1 (.DIODE(_06337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13219__A1 (.DIODE(_06337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13151__A1 (.DIODE(_06337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13083__A1 (.DIODE(_06337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12946__A1 (.DIODE(_06337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12878__A1 (.DIODE(_06337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12675__A1 (.DIODE(_06337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12597__A1 (.DIODE(_06337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13766__A1 (.DIODE(_06339_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13630__A1 (.DIODE(_06339_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13494__A1 (.DIODE(_06339_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13221__A1 (.DIODE(_06339_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13153__A1 (.DIODE(_06339_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13085__A1 (.DIODE(_06339_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12948__A1 (.DIODE(_06339_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12880__A1 (.DIODE(_06339_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12677__A1 (.DIODE(_06339_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12600__A1 (.DIODE(_06339_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13768__A1 (.DIODE(_06341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13632__A1 (.DIODE(_06341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13496__A1 (.DIODE(_06341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13223__A1 (.DIODE(_06341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13155__A1 (.DIODE(_06341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13087__A1 (.DIODE(_06341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12950__A1 (.DIODE(_06341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12882__A1 (.DIODE(_06341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12679__A1 (.DIODE(_06341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12603__A1 (.DIODE(_06341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13770__A1 (.DIODE(_06343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13634__A1 (.DIODE(_06343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13498__A1 (.DIODE(_06343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13225__A1 (.DIODE(_06343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13157__A1 (.DIODE(_06343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13089__A1 (.DIODE(_06343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12952__A1 (.DIODE(_06343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12884__A1 (.DIODE(_06343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12681__A1 (.DIODE(_06343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12606__A1 (.DIODE(_06343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13772__A1 (.DIODE(_06345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13636__A1 (.DIODE(_06345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13500__A1 (.DIODE(_06345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13227__A1 (.DIODE(_06345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13159__A1 (.DIODE(_06345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13091__A1 (.DIODE(_06345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12954__A1 (.DIODE(_06345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12886__A1 (.DIODE(_06345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12683__A1 (.DIODE(_06345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12609__A1 (.DIODE(_06345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13774__A1 (.DIODE(_06347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13638__A1 (.DIODE(_06347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13502__A1 (.DIODE(_06347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13229__A1 (.DIODE(_06347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13161__A1 (.DIODE(_06347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13093__A1 (.DIODE(_06347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12956__A1 (.DIODE(_06347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12888__A1 (.DIODE(_06347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12685__A1 (.DIODE(_06347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12612__A1 (.DIODE(_06347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13776__A1 (.DIODE(_06349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13640__A1 (.DIODE(_06349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13504__A1 (.DIODE(_06349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13231__A1 (.DIODE(_06349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13163__A1 (.DIODE(_06349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13095__A1 (.DIODE(_06349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12958__A1 (.DIODE(_06349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12890__A1 (.DIODE(_06349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12687__A1 (.DIODE(_06349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12615__A1 (.DIODE(_06349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13778__A1 (.DIODE(_06351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13642__A1 (.DIODE(_06351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13506__A1 (.DIODE(_06351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13233__A1 (.DIODE(_06351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13165__A1 (.DIODE(_06351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13097__A1 (.DIODE(_06351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12960__A1 (.DIODE(_06351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12892__A1 (.DIODE(_06351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12689__A1 (.DIODE(_06351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12618__A1 (.DIODE(_06351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13780__A1 (.DIODE(_06353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13644__A1 (.DIODE(_06353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13508__A1 (.DIODE(_06353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13235__A1 (.DIODE(_06353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13167__A1 (.DIODE(_06353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13099__A1 (.DIODE(_06353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12962__A1 (.DIODE(_06353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12894__A1 (.DIODE(_06353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12691__A1 (.DIODE(_06353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12621__A1 (.DIODE(_06353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13782__A1 (.DIODE(_06355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13646__A1 (.DIODE(_06355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13510__A1 (.DIODE(_06355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13237__A1 (.DIODE(_06355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13169__A1 (.DIODE(_06355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13101__A1 (.DIODE(_06355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12964__A1 (.DIODE(_06355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12896__A1 (.DIODE(_06355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12693__A1 (.DIODE(_06355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12624__A1 (.DIODE(_06355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12649__S (.DIODE(_06360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12647__S (.DIODE(_06360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12645__S (.DIODE(_06360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12643__S (.DIODE(_06360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12641__S (.DIODE(_06360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12639__S (.DIODE(_06360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12637__S (.DIODE(_06360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12635__S (.DIODE(_06360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12633__S (.DIODE(_06360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12631__S (.DIODE(_06360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12670__S (.DIODE(_06371_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12668__S (.DIODE(_06371_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12666__S (.DIODE(_06371_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12664__S (.DIODE(_06371_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12662__S (.DIODE(_06371_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12660__S (.DIODE(_06371_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12658__S (.DIODE(_06371_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12656__S (.DIODE(_06371_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12654__S (.DIODE(_06371_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12652__S (.DIODE(_06371_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12691__S (.DIODE(_06382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12689__S (.DIODE(_06382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12687__S (.DIODE(_06382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12685__S (.DIODE(_06382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12683__S (.DIODE(_06382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12681__S (.DIODE(_06382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12679__S (.DIODE(_06382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12677__S (.DIODE(_06382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12675__S (.DIODE(_06382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12673__S (.DIODE(_06382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12763__S (.DIODE(_06395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12761__S (.DIODE(_06395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12740__A (.DIODE(_06395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12719__A (.DIODE(_06395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12698__A (.DIODE(_06395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12717__S (.DIODE(_06396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12715__S (.DIODE(_06396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12713__S (.DIODE(_06396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12711__S (.DIODE(_06396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12709__S (.DIODE(_06396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12707__S (.DIODE(_06396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12705__S (.DIODE(_06396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12703__S (.DIODE(_06396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12701__S (.DIODE(_06396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12699__S (.DIODE(_06396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12738__S (.DIODE(_06407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12736__S (.DIODE(_06407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12734__S (.DIODE(_06407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12732__S (.DIODE(_06407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12730__S (.DIODE(_06407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12728__S (.DIODE(_06407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12726__S (.DIODE(_06407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12724__S (.DIODE(_06407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12722__S (.DIODE(_06407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12720__S (.DIODE(_06407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12759__S (.DIODE(_06418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12757__S (.DIODE(_06418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12755__S (.DIODE(_06418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12753__S (.DIODE(_06418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12751__S (.DIODE(_06418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12749__S (.DIODE(_06418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12747__S (.DIODE(_06418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12745__S (.DIODE(_06418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12743__S (.DIODE(_06418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12741__S (.DIODE(_06418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12803__A (.DIODE(_06440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12801__A (.DIODE(_06440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12799__A (.DIODE(_06440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12797__A (.DIODE(_06440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12795__A (.DIODE(_06440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12793__A (.DIODE(_06440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12791__A (.DIODE(_06440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12789__A (.DIODE(_06440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12787__A (.DIODE(_06440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12785__A (.DIODE(_06440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12824__A (.DIODE(_06451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12822__A (.DIODE(_06451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12820__A (.DIODE(_06451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12818__A (.DIODE(_06451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12816__A (.DIODE(_06451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12814__A (.DIODE(_06451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12812__A (.DIODE(_06451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12810__A (.DIODE(_06451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12808__A (.DIODE(_06451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12806__A (.DIODE(_06451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12852__S (.DIODE(_06466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12850__S (.DIODE(_06466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12848__S (.DIODE(_06466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12846__S (.DIODE(_06466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12844__S (.DIODE(_06466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12842__S (.DIODE(_06466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12840__S (.DIODE(_06466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12838__S (.DIODE(_06466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12836__S (.DIODE(_06466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12834__S (.DIODE(_06466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12873__S (.DIODE(_06477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12871__S (.DIODE(_06477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12869__S (.DIODE(_06477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12867__S (.DIODE(_06477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12865__S (.DIODE(_06477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12863__S (.DIODE(_06477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12861__S (.DIODE(_06477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12859__S (.DIODE(_06477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12857__S (.DIODE(_06477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12855__S (.DIODE(_06477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12894__S (.DIODE(_06488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12892__S (.DIODE(_06488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12890__S (.DIODE(_06488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12888__S (.DIODE(_06488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12886__S (.DIODE(_06488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12884__S (.DIODE(_06488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12882__S (.DIODE(_06488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12880__S (.DIODE(_06488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12878__S (.DIODE(_06488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12876__S (.DIODE(_06488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12966__S (.DIODE(_06501_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12964__S (.DIODE(_06501_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12943__A (.DIODE(_06501_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12922__A (.DIODE(_06501_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12901__A (.DIODE(_06501_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12920__S (.DIODE(_06502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12918__S (.DIODE(_06502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12916__S (.DIODE(_06502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12914__S (.DIODE(_06502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12912__S (.DIODE(_06502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12910__S (.DIODE(_06502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12908__S (.DIODE(_06502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12906__S (.DIODE(_06502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12904__S (.DIODE(_06502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12902__S (.DIODE(_06502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12941__S (.DIODE(_06513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12939__S (.DIODE(_06513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12937__S (.DIODE(_06513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12935__S (.DIODE(_06513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12933__S (.DIODE(_06513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12931__S (.DIODE(_06513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12929__S (.DIODE(_06513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12927__S (.DIODE(_06513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12925__S (.DIODE(_06513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12923__S (.DIODE(_06513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12962__S (.DIODE(_06524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12960__S (.DIODE(_06524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12958__S (.DIODE(_06524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12956__S (.DIODE(_06524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12954__S (.DIODE(_06524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12952__S (.DIODE(_06524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12950__S (.DIODE(_06524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12948__S (.DIODE(_06524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12946__S (.DIODE(_06524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12944__S (.DIODE(_06524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13035__S (.DIODE(_06538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13033__S (.DIODE(_06538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13012__A (.DIODE(_06538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12991__A (.DIODE(_06538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12970__A (.DIODE(_06538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12989__S (.DIODE(_06539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12987__S (.DIODE(_06539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12985__S (.DIODE(_06539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12983__S (.DIODE(_06539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12981__S (.DIODE(_06539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12979__S (.DIODE(_06539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12977__S (.DIODE(_06539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12975__S (.DIODE(_06539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12973__S (.DIODE(_06539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12971__S (.DIODE(_06539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13010__S (.DIODE(_06550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13008__S (.DIODE(_06550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13006__S (.DIODE(_06550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13004__S (.DIODE(_06550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13002__S (.DIODE(_06550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13000__S (.DIODE(_06550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12998__S (.DIODE(_06550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12996__S (.DIODE(_06550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12994__S (.DIODE(_06550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12992__S (.DIODE(_06550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13031__S (.DIODE(_06561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13029__S (.DIODE(_06561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13027__S (.DIODE(_06561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13025__S (.DIODE(_06561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13023__S (.DIODE(_06561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13021__S (.DIODE(_06561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13019__S (.DIODE(_06561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13017__S (.DIODE(_06561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13015__S (.DIODE(_06561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13013__S (.DIODE(_06561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13103__S (.DIODE(_06574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13101__S (.DIODE(_06574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13080__A (.DIODE(_06574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13059__A (.DIODE(_06574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13038__A (.DIODE(_06574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13057__S (.DIODE(_06575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13055__S (.DIODE(_06575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13053__S (.DIODE(_06575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13051__S (.DIODE(_06575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13049__S (.DIODE(_06575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13047__S (.DIODE(_06575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13045__S (.DIODE(_06575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13043__S (.DIODE(_06575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13041__S (.DIODE(_06575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13039__S (.DIODE(_06575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13078__S (.DIODE(_06586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13076__S (.DIODE(_06586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13074__S (.DIODE(_06586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13072__S (.DIODE(_06586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13070__S (.DIODE(_06586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13068__S (.DIODE(_06586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13066__S (.DIODE(_06586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13064__S (.DIODE(_06586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13062__S (.DIODE(_06586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13060__S (.DIODE(_06586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13099__S (.DIODE(_06597_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13097__S (.DIODE(_06597_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13095__S (.DIODE(_06597_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13093__S (.DIODE(_06597_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13091__S (.DIODE(_06597_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13089__S (.DIODE(_06597_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13087__S (.DIODE(_06597_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13085__S (.DIODE(_06597_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13083__S (.DIODE(_06597_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13081__S (.DIODE(_06597_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13171__S (.DIODE(_06610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13169__S (.DIODE(_06610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13148__A (.DIODE(_06610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13127__A (.DIODE(_06610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13106__A (.DIODE(_06610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13125__S (.DIODE(_06611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13123__S (.DIODE(_06611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13121__S (.DIODE(_06611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13119__S (.DIODE(_06611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13117__S (.DIODE(_06611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13115__S (.DIODE(_06611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13113__S (.DIODE(_06611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13111__S (.DIODE(_06611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13109__S (.DIODE(_06611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13107__S (.DIODE(_06611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13146__S (.DIODE(_06622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13144__S (.DIODE(_06622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13142__S (.DIODE(_06622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13140__S (.DIODE(_06622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13138__S (.DIODE(_06622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13136__S (.DIODE(_06622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13134__S (.DIODE(_06622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13132__S (.DIODE(_06622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13130__S (.DIODE(_06622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13128__S (.DIODE(_06622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13167__S (.DIODE(_06633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13165__S (.DIODE(_06633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13163__S (.DIODE(_06633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13161__S (.DIODE(_06633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13159__S (.DIODE(_06633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13157__S (.DIODE(_06633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13155__S (.DIODE(_06633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13153__S (.DIODE(_06633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13151__S (.DIODE(_06633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13149__S (.DIODE(_06633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13239__S (.DIODE(_06646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13237__S (.DIODE(_06646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13216__A (.DIODE(_06646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13195__A (.DIODE(_06646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13174__A (.DIODE(_06646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13193__S (.DIODE(_06647_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13191__S (.DIODE(_06647_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13189__S (.DIODE(_06647_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13187__S (.DIODE(_06647_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13185__S (.DIODE(_06647_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13183__S (.DIODE(_06647_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13181__S (.DIODE(_06647_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13179__S (.DIODE(_06647_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13177__S (.DIODE(_06647_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13175__S (.DIODE(_06647_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13214__S (.DIODE(_06658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13212__S (.DIODE(_06658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13210__S (.DIODE(_06658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13208__S (.DIODE(_06658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13206__S (.DIODE(_06658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13204__S (.DIODE(_06658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13202__S (.DIODE(_06658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13200__S (.DIODE(_06658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13198__S (.DIODE(_06658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13196__S (.DIODE(_06658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13235__S (.DIODE(_06669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13233__S (.DIODE(_06669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13231__S (.DIODE(_06669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13229__S (.DIODE(_06669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13227__S (.DIODE(_06669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13225__S (.DIODE(_06669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13223__S (.DIODE(_06669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13221__S (.DIODE(_06669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13219__S (.DIODE(_06669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13217__S (.DIODE(_06669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13308__S (.DIODE(_06683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13306__S (.DIODE(_06683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13285__A (.DIODE(_06683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13264__A (.DIODE(_06683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13243__A (.DIODE(_06683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13262__S (.DIODE(_06684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13260__S (.DIODE(_06684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13258__S (.DIODE(_06684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13256__S (.DIODE(_06684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13254__S (.DIODE(_06684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13252__S (.DIODE(_06684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13250__S (.DIODE(_06684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13248__S (.DIODE(_06684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13246__S (.DIODE(_06684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13244__S (.DIODE(_06684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13283__S (.DIODE(_06695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13281__S (.DIODE(_06695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13279__S (.DIODE(_06695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13277__S (.DIODE(_06695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13275__S (.DIODE(_06695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13273__S (.DIODE(_06695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13271__S (.DIODE(_06695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13269__S (.DIODE(_06695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13267__S (.DIODE(_06695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13265__S (.DIODE(_06695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13304__S (.DIODE(_06706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13302__S (.DIODE(_06706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13300__S (.DIODE(_06706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13298__S (.DIODE(_06706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13296__S (.DIODE(_06706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13294__S (.DIODE(_06706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13292__S (.DIODE(_06706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13290__S (.DIODE(_06706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13288__S (.DIODE(_06706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13286__S (.DIODE(_06706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13330__S (.DIODE(_06720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13328__S (.DIODE(_06720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13326__S (.DIODE(_06720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13324__S (.DIODE(_06720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13322__S (.DIODE(_06720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13320__S (.DIODE(_06720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13318__S (.DIODE(_06720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13316__S (.DIODE(_06720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13314__S (.DIODE(_06720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13312__S (.DIODE(_06720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13351__S (.DIODE(_06731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13349__S (.DIODE(_06731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13347__S (.DIODE(_06731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13345__S (.DIODE(_06731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13343__S (.DIODE(_06731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13341__S (.DIODE(_06731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13339__S (.DIODE(_06731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13337__S (.DIODE(_06731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13335__S (.DIODE(_06731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13333__S (.DIODE(_06731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13372__S (.DIODE(_06742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13370__S (.DIODE(_06742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13368__S (.DIODE(_06742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13366__S (.DIODE(_06742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13364__S (.DIODE(_06742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13362__S (.DIODE(_06742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13360__S (.DIODE(_06742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13358__S (.DIODE(_06742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13356__S (.DIODE(_06742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13354__S (.DIODE(_06742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13398__S (.DIODE(_06756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13396__S (.DIODE(_06756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13394__S (.DIODE(_06756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13392__S (.DIODE(_06756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13390__S (.DIODE(_06756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13388__S (.DIODE(_06756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13386__S (.DIODE(_06756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13384__S (.DIODE(_06756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13382__S (.DIODE(_06756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13380__S (.DIODE(_06756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13419__S (.DIODE(_06767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13417__S (.DIODE(_06767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13415__S (.DIODE(_06767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13413__S (.DIODE(_06767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13411__S (.DIODE(_06767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13409__S (.DIODE(_06767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13407__S (.DIODE(_06767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13405__S (.DIODE(_06767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13403__S (.DIODE(_06767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13401__S (.DIODE(_06767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13440__S (.DIODE(_06778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13438__S (.DIODE(_06778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13436__S (.DIODE(_06778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13434__S (.DIODE(_06778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13432__S (.DIODE(_06778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13430__S (.DIODE(_06778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13428__S (.DIODE(_06778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13426__S (.DIODE(_06778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13424__S (.DIODE(_06778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13422__S (.DIODE(_06778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13512__S (.DIODE(_06791_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13510__S (.DIODE(_06791_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13489__A (.DIODE(_06791_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13468__A (.DIODE(_06791_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13447__A (.DIODE(_06791_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13466__S (.DIODE(_06792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13464__S (.DIODE(_06792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13462__S (.DIODE(_06792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13460__S (.DIODE(_06792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13458__S (.DIODE(_06792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13456__S (.DIODE(_06792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13454__S (.DIODE(_06792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13452__S (.DIODE(_06792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13450__S (.DIODE(_06792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13448__S (.DIODE(_06792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13487__S (.DIODE(_06803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13485__S (.DIODE(_06803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13483__S (.DIODE(_06803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13481__S (.DIODE(_06803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13479__S (.DIODE(_06803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13477__S (.DIODE(_06803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13475__S (.DIODE(_06803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13473__S (.DIODE(_06803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13471__S (.DIODE(_06803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13469__S (.DIODE(_06803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13508__S (.DIODE(_06814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13506__S (.DIODE(_06814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13504__S (.DIODE(_06814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13502__S (.DIODE(_06814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13500__S (.DIODE(_06814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13498__S (.DIODE(_06814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13496__S (.DIODE(_06814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13494__S (.DIODE(_06814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13492__S (.DIODE(_06814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13490__S (.DIODE(_06814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13534__S (.DIODE(_06828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13532__S (.DIODE(_06828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13530__S (.DIODE(_06828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13528__S (.DIODE(_06828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13526__S (.DIODE(_06828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13524__S (.DIODE(_06828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13522__S (.DIODE(_06828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13520__S (.DIODE(_06828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13518__S (.DIODE(_06828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13516__S (.DIODE(_06828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13555__S (.DIODE(_06839_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13553__S (.DIODE(_06839_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13551__S (.DIODE(_06839_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13549__S (.DIODE(_06839_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13547__S (.DIODE(_06839_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13545__S (.DIODE(_06839_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13543__S (.DIODE(_06839_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13541__S (.DIODE(_06839_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13539__S (.DIODE(_06839_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13537__S (.DIODE(_06839_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13576__S (.DIODE(_06850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13574__S (.DIODE(_06850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13572__S (.DIODE(_06850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13570__S (.DIODE(_06850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13568__S (.DIODE(_06850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13566__S (.DIODE(_06850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13564__S (.DIODE(_06850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13562__S (.DIODE(_06850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13560__S (.DIODE(_06850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13558__S (.DIODE(_06850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13602__S (.DIODE(_06864_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13600__S (.DIODE(_06864_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13598__S (.DIODE(_06864_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13596__S (.DIODE(_06864_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13594__S (.DIODE(_06864_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13592__S (.DIODE(_06864_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13590__S (.DIODE(_06864_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13588__S (.DIODE(_06864_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13586__S (.DIODE(_06864_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13584__S (.DIODE(_06864_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13623__S (.DIODE(_06875_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13621__S (.DIODE(_06875_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13619__S (.DIODE(_06875_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13617__S (.DIODE(_06875_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13615__S (.DIODE(_06875_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13613__S (.DIODE(_06875_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13611__S (.DIODE(_06875_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13609__S (.DIODE(_06875_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13607__S (.DIODE(_06875_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13605__S (.DIODE(_06875_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13644__S (.DIODE(_06886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13642__S (.DIODE(_06886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13640__S (.DIODE(_06886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13638__S (.DIODE(_06886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13636__S (.DIODE(_06886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13634__S (.DIODE(_06886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13632__S (.DIODE(_06886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13630__S (.DIODE(_06886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13628__S (.DIODE(_06886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13626__S (.DIODE(_06886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13716__S (.DIODE(_06899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13714__S (.DIODE(_06899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13693__A (.DIODE(_06899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13672__A (.DIODE(_06899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13651__A (.DIODE(_06899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13670__S (.DIODE(_06900_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13668__S (.DIODE(_06900_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13666__S (.DIODE(_06900_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13664__S (.DIODE(_06900_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13662__S (.DIODE(_06900_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13660__S (.DIODE(_06900_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13658__S (.DIODE(_06900_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13656__S (.DIODE(_06900_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13654__S (.DIODE(_06900_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13652__S (.DIODE(_06900_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13691__S (.DIODE(_06911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13689__S (.DIODE(_06911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13687__S (.DIODE(_06911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13685__S (.DIODE(_06911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13683__S (.DIODE(_06911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13681__S (.DIODE(_06911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13679__S (.DIODE(_06911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13677__S (.DIODE(_06911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13675__S (.DIODE(_06911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13673__S (.DIODE(_06911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13712__S (.DIODE(_06922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13710__S (.DIODE(_06922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13708__S (.DIODE(_06922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13706__S (.DIODE(_06922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13704__S (.DIODE(_06922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13702__S (.DIODE(_06922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13700__S (.DIODE(_06922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13698__S (.DIODE(_06922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13696__S (.DIODE(_06922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13694__S (.DIODE(_06922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13738__S (.DIODE(_06936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13736__S (.DIODE(_06936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13734__S (.DIODE(_06936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13732__S (.DIODE(_06936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13730__S (.DIODE(_06936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13728__S (.DIODE(_06936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13726__S (.DIODE(_06936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13724__S (.DIODE(_06936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13722__S (.DIODE(_06936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13720__S (.DIODE(_06936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13759__S (.DIODE(_06947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13757__S (.DIODE(_06947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13755__S (.DIODE(_06947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13753__S (.DIODE(_06947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13751__S (.DIODE(_06947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13749__S (.DIODE(_06947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13747__S (.DIODE(_06947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13745__S (.DIODE(_06947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13743__S (.DIODE(_06947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13741__S (.DIODE(_06947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13780__S (.DIODE(_06958_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13778__S (.DIODE(_06958_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13776__S (.DIODE(_06958_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13774__S (.DIODE(_06958_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13772__S (.DIODE(_06958_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13770__S (.DIODE(_06958_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13768__S (.DIODE(_06958_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13766__S (.DIODE(_06958_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13764__S (.DIODE(_06958_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13762__S (.DIODE(_06958_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13802__A (.DIODE(_06971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13801__A (.DIODE(_06971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13800__A (.DIODE(_06971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13799__A (.DIODE(_06971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13798__A (.DIODE(_06971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13797__A (.DIODE(_06971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13796__A (.DIODE(_06971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13795__A (.DIODE(_06971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13794__A (.DIODE(_06971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13793__A (.DIODE(_06971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13813__A (.DIODE(_06972_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13812__A (.DIODE(_06972_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13811__A (.DIODE(_06972_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13810__A (.DIODE(_06972_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13809__A (.DIODE(_06972_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13808__A (.DIODE(_06972_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13807__A (.DIODE(_06972_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13806__A (.DIODE(_06972_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13805__A (.DIODE(_06972_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13804__A (.DIODE(_06972_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13824__A (.DIODE(_06973_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13823__A (.DIODE(_06973_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13822__A (.DIODE(_06973_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13821__A (.DIODE(_06973_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13820__A (.DIODE(_06973_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13819__A (.DIODE(_06973_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13818__A (.DIODE(_06973_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13817__A (.DIODE(_06973_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13816__A (.DIODE(_06973_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13815__A (.DIODE(_06973_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13868__A (.DIODE(_06977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13867__A (.DIODE(_06977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13866__A (.DIODE(_06977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13865__A (.DIODE(_06977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13864__A (.DIODE(_06977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13863__A (.DIODE(_06977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13862__A (.DIODE(_06977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13861__A (.DIODE(_06977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13860__A (.DIODE(_06977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13859__A (.DIODE(_06977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13991__A (.DIODE(_06980_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13980__A (.DIODE(_06980_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13969__A (.DIODE(_06980_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13958__A (.DIODE(_06980_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13947__A (.DIODE(_06980_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13936__A (.DIODE(_06980_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13925__A (.DIODE(_06980_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13914__A (.DIODE(_06980_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13903__A (.DIODE(_06980_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13892__A (.DIODE(_06980_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13902__A (.DIODE(_06981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13901__A (.DIODE(_06981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13900__A (.DIODE(_06981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13899__A (.DIODE(_06981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13898__A (.DIODE(_06981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13897__A (.DIODE(_06981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13896__A (.DIODE(_06981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13895__A (.DIODE(_06981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13894__A (.DIODE(_06981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13893__A (.DIODE(_06981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13924__A (.DIODE(_06983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13923__A (.DIODE(_06983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13922__A (.DIODE(_06983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13921__A (.DIODE(_06983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13920__A (.DIODE(_06983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13919__A (.DIODE(_06983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13918__A (.DIODE(_06983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13917__A (.DIODE(_06983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13916__A (.DIODE(_06983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13915__A (.DIODE(_06983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13935__A (.DIODE(_06984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13934__A (.DIODE(_06984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13933__A (.DIODE(_06984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13932__A (.DIODE(_06984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13931__A (.DIODE(_06984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13930__A (.DIODE(_06984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13929__A (.DIODE(_06984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13928__A (.DIODE(_06984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13927__A (.DIODE(_06984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13926__A (.DIODE(_06984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13990__A (.DIODE(_06989_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13989__A (.DIODE(_06989_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13988__A (.DIODE(_06989_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13987__A (.DIODE(_06989_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13986__A (.DIODE(_06989_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13985__A (.DIODE(_06989_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13984__A (.DIODE(_06989_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13983__A (.DIODE(_06989_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13982__A (.DIODE(_06989_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13981__A (.DIODE(_06989_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14001__A (.DIODE(_06990_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14000__A (.DIODE(_06990_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13999__A (.DIODE(_06990_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13998__A (.DIODE(_06990_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13997__A (.DIODE(_06990_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13996__A (.DIODE(_06990_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13995__A (.DIODE(_06990_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13994__A (.DIODE(_06990_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13993__A (.DIODE(_06990_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13992__A (.DIODE(_06990_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14012__A (.DIODE(_06991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14011__A (.DIODE(_06991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14010__A (.DIODE(_06991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14009__A (.DIODE(_06991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14008__A (.DIODE(_06991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14007__A (.DIODE(_06991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14006__A (.DIODE(_06991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14005__A (.DIODE(_06991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14004__A (.DIODE(_06991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14003__A (.DIODE(_06991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14023__A (.DIODE(_06992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14022__A (.DIODE(_06992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14021__A (.DIODE(_06992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14020__A (.DIODE(_06992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14019__A (.DIODE(_06992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14018__A (.DIODE(_06992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14017__A (.DIODE(_06992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14016__A (.DIODE(_06992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14015__A (.DIODE(_06992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14014__A (.DIODE(_06992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14102__A (.DIODE(_06993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14101__A (.DIODE(_06993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14032__A (.DIODE(_06993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14031__A (.DIODE(_06993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14030__A (.DIODE(_06993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14029__A (.DIODE(_06993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14028__A (.DIODE(_06993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14027__A (.DIODE(_06993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14026__A (.DIODE(_06993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14025__A (.DIODE(_06993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14053__S (.DIODE(_06995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14051__S (.DIODE(_06995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14049__S (.DIODE(_06995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14047__S (.DIODE(_06995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14045__S (.DIODE(_06995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14043__S (.DIODE(_06995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14041__S (.DIODE(_06995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14039__S (.DIODE(_06995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14037__S (.DIODE(_06995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14035__S (.DIODE(_06995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14074__S (.DIODE(_07006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14072__S (.DIODE(_07006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14070__S (.DIODE(_07006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14068__S (.DIODE(_07006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14066__S (.DIODE(_07006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14064__S (.DIODE(_07006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14062__S (.DIODE(_07006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14060__S (.DIODE(_07006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14058__S (.DIODE(_07006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14056__S (.DIODE(_07006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14095__S (.DIODE(_07017_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14093__S (.DIODE(_07017_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14091__S (.DIODE(_07017_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14089__S (.DIODE(_07017_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14087__S (.DIODE(_07017_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14085__S (.DIODE(_07017_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14083__S (.DIODE(_07017_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14081__S (.DIODE(_07017_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14079__S (.DIODE(_07017_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14077__S (.DIODE(_07017_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14113__A (.DIODE(_07030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14112__A (.DIODE(_07030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14111__A (.DIODE(_07030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14110__A (.DIODE(_07030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14109__A (.DIODE(_07030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14108__A (.DIODE(_07030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14107__A (.DIODE(_07030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14106__A (.DIODE(_07030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14105__A (.DIODE(_07030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14104__A (.DIODE(_07030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14124__A (.DIODE(_07031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14123__A (.DIODE(_07031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14122__A (.DIODE(_07031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14121__A (.DIODE(_07031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14120__A (.DIODE(_07031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14119__A (.DIODE(_07031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14118__A (.DIODE(_07031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14117__A (.DIODE(_07031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14116__A (.DIODE(_07031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14115__A (.DIODE(_07031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10529__A (.DIODE(\barrel_shifter_right.arith ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10290__A0 (.DIODE(\barrel_shifter_right.arith ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07385__A (.DIODE(\barrel_shifter_right.arith ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07108__A (.DIODE(\barrel_shifter_right.arith ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07107__B (.DIODE(\barrel_shifter_right.arith ));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_A (.DIODE(clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__10177__A_N (.DIODE(\instr[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09738__A (.DIODE(\instr[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07880__A0 (.DIODE(\instr[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07521__A (.DIODE(\instr[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07509__A (.DIODE(\instr[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07499__A1 (.DIODE(\instr[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07498__A (.DIODE(\instr[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07367__A (.DIODE(\instr[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07359__A_N (.DIODE(\instr[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07039__A (.DIODE(\instr[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10477__A0 (.DIODE(\leorv32_alu.input1[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09760__A2 (.DIODE(\leorv32_alu.input1[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07409__B (.DIODE(\leorv32_alu.input1[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07313__A (.DIODE(\leorv32_alu.input1[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07282__A (.DIODE(\leorv32_alu.input1[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11401__A1 (.DIODE(\leorv32_alu.input1[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11368__A1 (.DIODE(\leorv32_alu.input1[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10491__A1 (.DIODE(\leorv32_alu.input1[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10472__A0 (.DIODE(\leorv32_alu.input1[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10374__A1 (.DIODE(\leorv32_alu.input1[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08259__A0 (.DIODE(\leorv32_alu.input1[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07371__B (.DIODE(\leorv32_alu.input1[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07370__B (.DIODE(\leorv32_alu.input1[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07369__B (.DIODE(\leorv32_alu.input1[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07221__A (.DIODE(\leorv32_alu.input1[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10459__A1 (.DIODE(\leorv32_alu.input1[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10357__A (.DIODE(\leorv32_alu.input1[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10355__A (.DIODE(\leorv32_alu.input1[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08236__A1 (.DIODE(\leorv32_alu.input1[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07457__B (.DIODE(\leorv32_alu.input1[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07369__A (.DIODE(\leorv32_alu.input1[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07220__A (.DIODE(\leorv32_alu.input1[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11427__A (.DIODE(\leorv32_alu.input1[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10568__D (.DIODE(\leorv32_alu.input1[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10512__A1 (.DIODE(\leorv32_alu.input1[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10448__A0 (.DIODE(\leorv32_alu.input1[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10347__A (.DIODE(\leorv32_alu.input1[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08213__A1 (.DIODE(\leorv32_alu.input1[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07469__B (.DIODE(\leorv32_alu.input1[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07459__B (.DIODE(\leorv32_alu.input1[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07368__B (.DIODE(\leorv32_alu.input1[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07218__A (.DIODE(\leorv32_alu.input1[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11422__A (.DIODE(\leorv32_alu.input1[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11421__A (.DIODE(\leorv32_alu.input1[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10568__C (.DIODE(\leorv32_alu.input1[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10480__A1 (.DIODE(\leorv32_alu.input1[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08189__A1 (.DIODE(\leorv32_alu.input1[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07461__B (.DIODE(\leorv32_alu.input1[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07217__A (.DIODE(\leorv32_alu.input1[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10568__B (.DIODE(\leorv32_alu.input1[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10497__A1 (.DIODE(\leorv32_alu.input1[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10479__A0 (.DIODE(\leorv32_alu.input1[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10384__A (.DIODE(\leorv32_alu.input1[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10383__A (.DIODE(\leorv32_alu.input1[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08167__A1 (.DIODE(\leorv32_alu.input1[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07239__A1 (.DIODE(\leorv32_alu.input1[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07209__A (.DIODE(\leorv32_alu.input1[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10568__A (.DIODE(\leorv32_alu.input1[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10511__A0 (.DIODE(\leorv32_alu.input1[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10449__A1 (.DIODE(\leorv32_alu.input1[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10380__A (.DIODE(\leorv32_alu.input1[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10379__A (.DIODE(\leorv32_alu.input1[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08136__A1 (.DIODE(\leorv32_alu.input1[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07208__A (.DIODE(\leorv32_alu.input1[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11571__A1 (.DIODE(\leorv32_alu.input1[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11534__A1 (.DIODE(\leorv32_alu.input1[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10569__D (.DIODE(\leorv32_alu.input1[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10517__A1 (.DIODE(\leorv32_alu.input1[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10458__A0 (.DIODE(\leorv32_alu.input1[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10421__A1 (.DIODE(\leorv32_alu.input1[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10420__A1 (.DIODE(\leorv32_alu.input1[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08109__A1 (.DIODE(\leorv32_alu.input1[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07214__B2 (.DIODE(\leorv32_alu.input1[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07211__A (.DIODE(\leorv32_alu.input1[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11570__A (.DIODE(\leorv32_alu.input1[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10569__C (.DIODE(\leorv32_alu.input1[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10490__A0 (.DIODE(\leorv32_alu.input1[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10473__A1 (.DIODE(\leorv32_alu.input1[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10392__A (.DIODE(\leorv32_alu.input1[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10391__A (.DIODE(\leorv32_alu.input1[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08084__A1 (.DIODE(\leorv32_alu.input1[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07206__A (.DIODE(\leorv32_alu.input1[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11586__A (.DIODE(\leorv32_alu.input1[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11585__A (.DIODE(\leorv32_alu.input1[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10569__A (.DIODE(\leorv32_alu.input1[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10520__A0 (.DIODE(\leorv32_alu.input1[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10456__A1 (.DIODE(\leorv32_alu.input1[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10400__A (.DIODE(\leorv32_alu.input1[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10399__A (.DIODE(\leorv32_alu.input1[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08036__A1 (.DIODE(\leorv32_alu.input1[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07205__A1 (.DIODE(\leorv32_alu.input1[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07203__B2 (.DIODE(\leorv32_alu.input1[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11643__A1 (.DIODE(\leorv32_alu.input1[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10570__B (.DIODE(\leorv32_alu.input1[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10509__A1 (.DIODE(\leorv32_alu.input1[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10441__A0 (.DIODE(\leorv32_alu.input1[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10425__A1 (.DIODE(\leorv32_alu.input1[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10410__A (.DIODE(\leorv32_alu.input1[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07998__A0 (.DIODE(\leorv32_alu.input1[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07311__A (.DIODE(\leorv32_alu.input1[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07203__A1 (.DIODE(\leorv32_alu.input1[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07200__A (.DIODE(\leorv32_alu.input1[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11648__A2 (.DIODE(\leorv32_alu.input1[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10570__A (.DIODE(\leorv32_alu.input1[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10500__A0 (.DIODE(\leorv32_alu.input1[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10477__A1 (.DIODE(\leorv32_alu.input1[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10426__A (.DIODE(\leorv32_alu.input1[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10403__A (.DIODE(\leorv32_alu.input1[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07963__A1 (.DIODE(\leorv32_alu.input1[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07201__B (.DIODE(\leorv32_alu.input1[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07197__A_N (.DIODE(\leorv32_alu.input1[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10804__A (.DIODE(\leorv32_alu.input1[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10803__A (.DIODE(\leorv32_alu.input1[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10565__C (.DIODE(\leorv32_alu.input1[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10517__A0 (.DIODE(\leorv32_alu.input1[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10458__A1 (.DIODE(\leorv32_alu.input1[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08604__A0 (.DIODE(\leorv32_alu.input1[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07417__B (.DIODE(\leorv32_alu.input1[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07397__B (.DIODE(\leorv32_alu.input1[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07269__A (.DIODE(\leorv32_alu.input1[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10837__A1_N (.DIODE(\leorv32_alu.input1[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10835__A (.DIODE(\leorv32_alu.input1[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10565__B (.DIODE(\leorv32_alu.input1[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10511__A1 (.DIODE(\leorv32_alu.input1[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10449__A0 (.DIODE(\leorv32_alu.input1[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07420__B (.DIODE(\leorv32_alu.input1[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07395__B (.DIODE(\leorv32_alu.input1[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07294__B2 (.DIODE(\leorv32_alu.input1[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07293__B1 (.DIODE(\leorv32_alu.input1[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07273__A (.DIODE(\leorv32_alu.input1[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10567__D (.DIODE(\leorv32_alu.input1[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10480__A0 (.DIODE(\leorv32_alu.input1[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10300__A (.DIODE(\leorv32_alu.input1[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10299__A (.DIODE(\leorv32_alu.input1[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08534__A0 (.DIODE(\leorv32_alu.input1[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07425__B (.DIODE(\leorv32_alu.input1[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07424__B (.DIODE(\leorv32_alu.input1[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07260__A (.DIODE(\leorv32_alu.input1[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(mem_rbusy));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(mem_rdata[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(mem_rdata[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_A (.DIODE(mem_rdata[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_A (.DIODE(mem_rdata[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_A (.DIODE(mem_rdata[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_A (.DIODE(mem_rdata[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_A (.DIODE(mem_rdata[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_A (.DIODE(mem_rdata[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_A (.DIODE(mem_rdata[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_A (.DIODE(mem_rdata[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_A (.DIODE(mem_rdata[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_A (.DIODE(mem_rdata[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_A (.DIODE(mem_rdata[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_A (.DIODE(mem_rdata[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_A (.DIODE(mem_rdata[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_A (.DIODE(mem_rdata[23]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_A (.DIODE(mem_rdata[24]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_A (.DIODE(mem_rdata[25]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_A (.DIODE(mem_rdata[26]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_A (.DIODE(mem_rdata[27]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_A (.DIODE(mem_rdata[28]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_A (.DIODE(mem_rdata[29]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_A (.DIODE(mem_rdata[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input25_A (.DIODE(mem_rdata[30]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input26_A (.DIODE(mem_rdata[31]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input27_A (.DIODE(mem_rdata[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input28_A (.DIODE(mem_rdata[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input29_A (.DIODE(mem_rdata[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input30_A (.DIODE(mem_rdata[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input31_A (.DIODE(mem_rdata[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input32_A (.DIODE(mem_rdata[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input33_A (.DIODE(mem_rdata[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input34_A (.DIODE(mem_wbusy));
 sky130_fd_sc_hd__diode_2 ANTENNA_input35_A (.DIODE(mhartid_0));
 sky130_fd_sc_hd__diode_2 ANTENNA__12806__B (.DIODE(\regs[0][19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09272__A0 (.DIODE(\regs[0][19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08265__A0 (.DIODE(\regs[0][19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12759__A1 (.DIODE(\regs[4][29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09033__A0 (.DIODE(\regs[4][29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08005__A0 (.DIODE(\regs[4][29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_input36_A (.DIODE(reset));
 sky130_fd_sc_hd__diode_2 ANTENNA__10615__A0 (.DIODE(\rs2_content[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10236__A1 (.DIODE(\rs2_content[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09976__B2 (.DIODE(\rs2_content[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09952__B2 (.DIODE(\rs2_content[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09926__B2 (.DIODE(\rs2_content[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09910__A (.DIODE(\rs2_content[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09719__A1 (.DIODE(\rs2_content[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07315__A2 (.DIODE(\rs2_content[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07312__A (.DIODE(\rs2_content[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07283__B1 (.DIODE(\rs2_content[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10290__A1 (.DIODE(\rs2_content[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09985__A1 (.DIODE(\rs2_content[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09932__A1 (.DIODE(\rs2_content[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09492__A0 (.DIODE(\rs2_content[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07256__A (.DIODE(\rs2_content[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11038__A1 (.DIODE(\rs2_content[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10293__A1 (.DIODE(\rs2_content[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09988__A1 (.DIODE(\rs2_content[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09935__A1 (.DIODE(\rs2_content[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09469__A1 (.DIODE(\rs2_content[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07254__A (.DIODE(\rs2_content[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10284__A1 (.DIODE(\rs2_content[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10283__A1 (.DIODE(\rs2_content[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09992__A1 (.DIODE(\rs2_content[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09939__A1 (.DIODE(\rs2_content[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09447__A1 (.DIODE(\rs2_content[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07251__A (.DIODE(\rs2_content[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10279__A1 (.DIODE(\rs2_content[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09996__A1 (.DIODE(\rs2_content[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09942__A1 (.DIODE(\rs2_content[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09425__A1 (.DIODE(\rs2_content[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07250__A (.DIODE(\rs2_content[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10273__A (.DIODE(\rs2_content[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10000__A1 (.DIODE(\rs2_content[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09945__A1 (.DIODE(\rs2_content[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09402__A1 (.DIODE(\rs2_content[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07248__A (.DIODE(\rs2_content[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10270__A1 (.DIODE(\rs2_content[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10004__A1 (.DIODE(\rs2_content[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09948__A1 (.DIODE(\rs2_content[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07247__A (.DIODE(\rs2_content[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10341__A1 (.DIODE(\rs2_content[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10339__A1 (.DIODE(\rs2_content[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09952__A1 (.DIODE(\rs2_content[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09357__A1 (.DIODE(\rs2_content[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07306__A1_N (.DIODE(\rs2_content[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07228__B_N (.DIODE(\rs2_content[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10334__A1 (.DIODE(\rs2_content[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09955__A1 (.DIODE(\rs2_content[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09335__A1 (.DIODE(\rs2_content[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07230__A_N (.DIODE(\rs2_content[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07227__B_N (.DIODE(\rs2_content[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10322__A1 (.DIODE(\rs2_content[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09958__A1 (.DIODE(\rs2_content[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09312__A0 (.DIODE(\rs2_content[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07225__A (.DIODE(\rs2_content[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10327__A1 (.DIODE(\rs2_content[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09961__A1 (.DIODE(\rs2_content[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09289__A1 (.DIODE(\rs2_content[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07224__A (.DIODE(\rs2_content[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10438__A0 (.DIODE(\rs2_content[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10232__A (.DIODE(\rs2_content[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09980__B2 (.DIODE(\rs2_content[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09955__B2 (.DIODE(\rs2_content[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09929__B2 (.DIODE(\rs2_content[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09912__A (.DIODE(\rs2_content[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07285__A (.DIODE(\rs2_content[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07283__A2 (.DIODE(\rs2_content[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10354__A1 (.DIODE(\rs2_content[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09967__A1 (.DIODE(\rs2_content[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09244__A1 (.DIODE(\rs2_content[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07235__B (.DIODE(\rs2_content[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07222__A2 (.DIODE(\rs2_content[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10382__A1 (.DIODE(\rs2_content[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09976__A1 (.DIODE(\rs2_content[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09167__A1 (.DIODE(\rs2_content[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07237__A (.DIODE(\rs2_content[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07210__B1 (.DIODE(\rs2_content[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10378__A1 (.DIODE(\rs2_content[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09980__A1 (.DIODE(\rs2_content[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09139__A0 (.DIODE(\rs2_content[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07212__B1 (.DIODE(\rs2_content[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07210__A2 (.DIODE(\rs2_content[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10390__A1 (.DIODE(\rs2_content[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09987__A1 (.DIODE(\rs2_content[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09093__A1 (.DIODE(\rs2_content[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07214__A2_N (.DIODE(\rs2_content[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07207__B (.DIODE(\rs2_content[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10405__A1 (.DIODE(\rs2_content[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09991__A1 (.DIODE(\rs2_content[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09068__A0 (.DIODE(\rs2_content[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07204__A (.DIODE(\rs2_content[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11584__A1 (.DIODE(\rs2_content[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10398__A1 (.DIODE(\rs2_content[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09995__A1 (.DIODE(\rs2_content[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07199__A (.DIODE(\rs2_content[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10411__A1 (.DIODE(\rs2_content[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10409__A1 (.DIODE(\rs2_content[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09999__A1 (.DIODE(\rs2_content[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08993__A1 (.DIODE(\rs2_content[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07202__A2 (.DIODE(\rs2_content[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07198__A (.DIODE(\rs2_content[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10402__A1 (.DIODE(\rs2_content[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10003__A1 (.DIODE(\rs2_content[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08945__A1 (.DIODE(\rs2_content[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07201__A_N (.DIODE(\rs2_content[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07197__B (.DIODE(\rs2_content[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10444__A0 (.DIODE(\rs2_content[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10253__A1 (.DIODE(\rs2_content[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09991__B2 (.DIODE(\rs2_content[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09964__B2 (.DIODE(\rs2_content[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09939__B2 (.DIODE(\rs2_content[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09918__A (.DIODE(\rs2_content[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09628__A1 (.DIODE(\rs2_content[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07317__A2 (.DIODE(\rs2_content[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07289__A2 (.DIODE(\rs2_content[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07275__B1 (.DIODE(\rs2_content[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10224__A1 (.DIODE(\rs2_content[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09995__B2 (.DIODE(\rs2_content[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09967__B2 (.DIODE(\rs2_content[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09942__B2 (.DIODE(\rs2_content[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09920__A (.DIODE(\rs2_content[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09606__A1 (.DIODE(\rs2_content[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07293__A1_N (.DIODE(\rs2_content[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07275__A2 (.DIODE(\rs2_content[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10262__A1 (.DIODE(\rs2_content[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09999__B2 (.DIODE(\rs2_content[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09970__B2 (.DIODE(\rs2_content[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09945__B2 (.DIODE(\rs2_content[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09922__A (.DIODE(\rs2_content[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09583__A1 (.DIODE(\rs2_content[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07292__A (.DIODE(\rs2_content[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07274__B1 (.DIODE(\rs2_content[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10221__A1 (.DIODE(\rs2_content[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10003__B2 (.DIODE(\rs2_content[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09973__B2 (.DIODE(\rs2_content[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09948__B2 (.DIODE(\rs2_content[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09924__A (.DIODE(\rs2_content[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09561__A1 (.DIODE(\rs2_content[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07316__A2 (.DIODE(\rs2_content[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07291__A (.DIODE(\rs2_content[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07274__A2 (.DIODE(\rs2_content[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10298__A1 (.DIODE(\rs2_content[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09977__A1 (.DIODE(\rs2_content[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09926__A1 (.DIODE(\rs2_content[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09538__A0 (.DIODE(\rs2_content[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07296__B (.DIODE(\rs2_content[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07261__A1_N (.DIODE(\rs2_content[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10303__A1 (.DIODE(\rs2_content[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09981__A1 (.DIODE(\rs2_content[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09929__A1 (.DIODE(\rs2_content[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09515__A1 (.DIODE(\rs2_content[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07257__A (.DIODE(\rs2_content[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09732__A1 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__09730__A1 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__08718__A (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07779__A (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__10557__A1 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__10556__A1 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__07887__A1 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__11012__A1 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__10640__A0 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__07866__A1 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__11050__A1 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__10681__A0 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__07863__A1 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__11056__A1 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__10768__A0 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__07860__A1 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__11096__A1 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__10777__A0 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__07857__A1 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__11130__A1 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__10818__A0 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__07855__A1 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__11228__A (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__10862__A0 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__07909__A (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__07893__A (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__07846__A (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__07991__A (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__07964__A (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__07947__A (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__07928__A (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__07903__A (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__07896__A (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__07841__A (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__11237__A1 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__10595__B2 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__08589__C1 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__08519__C1 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__08361__C1 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__07976__A (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__07919__A (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__07890__A (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__07836__A (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__11285__A1 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__10642__B2 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__08031__A (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__07922__A (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__07831__A (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__11291__A1 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__10683__B2 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__08602__B1 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__08532__B1 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__08374__B1 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__07995__A (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__07960__A (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__07826__A (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__10595__A1 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__07885__A1 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__09061__A (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__08927__A (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__08895__A (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__07820__A (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__09639__S1 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__09526__S1 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__09062__A (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__08930__A (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__08908__A (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__08903__A (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__08897__A (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__07815__A (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__11407__A1 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__10820__B2 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__09636__C1 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__09523__C1 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__09477__C1 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__09297__C1 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__08912__A (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__08901__A (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__08892__A (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__07809__A (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__11438__A1 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__08924__A (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__08915__A (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__07804__A (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__11475__A1 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__10553__A1 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__09649__B1 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__09536__B1 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__09490__B1 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__09310__B1 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__09188__B1 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__09137__B1 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__08891__A (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__07799__A (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__11500__A1 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__10593__A1 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__07797__A1 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__11525__A1 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__10640__A1 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__07795__A1 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__11549__A1 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__10681__A1 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__07793__A1 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__11578__A1 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__10768__A1 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__07791__A1 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__11606__A1 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__10777__A1 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__07789__A1 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__10642__A1 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__07883__A1 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__11632__A1 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__10818__A1 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__07787__A1 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__11657__A1 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__10862__A1 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__07785__A1 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__10683__A1 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__07880__A1 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__10770__A1 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__07878__A1 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__10779__A1 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__07876__A1 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__10820__A1 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__07874__A1 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__10866__A1 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__10860__A1 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__07872__A1 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__10909__A1 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__10553__A0 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__07870__A1 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__10950__A1 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__10593__A0 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__07868__A1 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__09730__A2 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__08718__B (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__10215__D_N (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA_output37_A (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_output53_A (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA_output55_A (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA_output56_A (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA_output76_A (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_output77_A (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_output78_A (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_output79_A (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_output80_A (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA_output81_A (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA_output82_A (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_output83_A (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA_output85_A (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_output86_A (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA_output94_A (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__09924__B (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__09922__B (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__09920__B (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__09918__B (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__09916__B (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__09914__B (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__09912__B (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__09910__B (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA_output95_A (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA_output96_A (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_output97_A (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_1_0_clk_A (.DIODE(clknet_1_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_0_0_clk_A (.DIODE(clknet_1_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_3_0_clk_A (.DIODE(clknet_1_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_2_0_clk_A (.DIODE(clknet_1_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_1_0_clk_A (.DIODE(clknet_2_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_0_0_clk_A (.DIODE(clknet_2_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_3_0_clk_A (.DIODE(clknet_2_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_2_0_clk_A (.DIODE(clknet_2_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_5_0_clk_A (.DIODE(clknet_2_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_4_0_clk_A (.DIODE(clknet_2_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_7_0_clk_A (.DIODE(clknet_2_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_6_0_clk_A (.DIODE(clknet_2_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_1_0_clk_A (.DIODE(clknet_3_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_0_0_clk_A (.DIODE(clknet_3_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_3_0_clk_A (.DIODE(clknet_3_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_2_0_clk_A (.DIODE(clknet_3_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_5_0_clk_A (.DIODE(clknet_3_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_4_0_clk_A (.DIODE(clknet_3_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_7_0_clk_A (.DIODE(clknet_3_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_6_0_clk_A (.DIODE(clknet_3_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_11_0_clk_A (.DIODE(clknet_3_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_10_0_clk_A (.DIODE(clknet_3_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_13_0_clk_A (.DIODE(clknet_3_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_12_0_clk_A (.DIODE(clknet_3_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_15_0_clk_A (.DIODE(clknet_3_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_14_0_clk_A (.DIODE(clknet_3_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_135_clk_A (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_134_clk_A (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_133_clk_A (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_132_clk_A (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_131_clk_A (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_130_clk_A (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_129_clk_A (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_2_clk_A (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_1_clk_A (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_0_clk_A (.DIODE(clknet_4_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_128_clk_A (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_127_clk_A (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_126_clk_A (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_125_clk_A (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_124_clk_A (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_123_clk_A (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_122_clk_A (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_109_clk_A (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_108_clk_A (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_107_clk_A (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_106_clk_A (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_105_clk_A (.DIODE(clknet_4_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_121_clk_A (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_14_clk_A (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_13_clk_A (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_12_clk_A (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_7_clk_A (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_6_clk_A (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_5_clk_A (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_4_clk_A (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_3_clk_A (.DIODE(clknet_4_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_120_clk_A (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_119_clk_A (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_118_clk_A (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_117_clk_A (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_116_clk_A (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_114_clk_A (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_15_clk_A (.DIODE(clknet_4_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_opt_1_0_clk_A (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_111_clk_A (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_110_clk_A (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_104_clk_A (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_103_clk_A (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_102_clk_A (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_101_clk_A (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_100_clk_A (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_99_clk_A (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_98_clk_A (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_97_clk_A (.DIODE(clknet_4_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_96_clk_A (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_95_clk_A (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_94_clk_A (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_93_clk_A (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_92_clk_A (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_91_clk_A (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_90_clk_A (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_88_clk_A (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_87_clk_A (.DIODE(clknet_4_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_115_clk_A (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_112_clk_A (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_78_clk_A (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_77_clk_A (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_76_clk_A (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_75_clk_A (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_74_clk_A (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_73_clk_A (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_72_clk_A (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_70_clk_A (.DIODE(clknet_4_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_89_clk_A (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_86_clk_A (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_85_clk_A (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_84_clk_A (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_83_clk_A (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_82_clk_A (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_81_clk_A (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_80_clk_A (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_79_clk_A (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_65_clk_A (.DIODE(clknet_4_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_30_clk_A (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_29_clk_A (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_28_clk_A (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_27_clk_A (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_25_clk_A (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_10_clk_A (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_9_clk_A (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_8_clk_A (.DIODE(clknet_4_8_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_26_clk_A (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_24_clk_A (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_23_clk_A (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_22_clk_A (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_21_clk_A (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_20_clk_A (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_17_clk_A (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_16_clk_A (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_11_clk_A (.DIODE(clknet_4_9_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_38_clk_A (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_37_clk_A (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_36_clk_A (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_35_clk_A (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_34_clk_A (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_33_clk_A (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_32_clk_A (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_31_clk_A (.DIODE(clknet_4_10_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_50_clk_A (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_49_clk_A (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_opt_2_0_clk_A (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_44_clk_A (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_43_clk_A (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_42_clk_A (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_41_clk_A (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_40_clk_A (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_39_clk_A (.DIODE(clknet_4_11_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_71_clk_A (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__15249__CLK (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_56_clk_A (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_55_clk_A (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_54_clk_A (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_19_clk_A (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_opt_3_0_clk_A (.DIODE(clknet_4_12_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_69_clk_A (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_68_clk_A (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_67_clk_A (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_66_clk_A (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_64_clk_A (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_63_clk_A (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_62_clk_A (.DIODE(clknet_4_13_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_57_clk_A (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_53_clk_A (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_52_clk_A (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_51_clk_A (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_48_clk_A (.DIODE(clknet_4_14_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_61_clk_A (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_60_clk_A (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_59_clk_A (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_47_clk_A (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_46_clk_A (.DIODE(clknet_4_15_0_clk));
 sky130_fd_sc_hd__decap_3 FILLER_0_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_482 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_632 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_795 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_977 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_990 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1002 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1057 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_470 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_535 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_646 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_715 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_758 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_831 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_984 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_996 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1052 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1058 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_235 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_599 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_672 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_731 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_803 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_859 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_873 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_879 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_891 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_488 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_547 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_772 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_831 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_887 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_266 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_332 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_438 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_574 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_593 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_744 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_803 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_859 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_891 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1057 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_303 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_528 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_565 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_646 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_702 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_831 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_887 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_901 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_913 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_202 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_263 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_288 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_661 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_788 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_800 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_859 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_903 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1052 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1058 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_292 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_386 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_526 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_548 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_640 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_646 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_691 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_831 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_887 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_913 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_919 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_931 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_226 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_576 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_627 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_663 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_676 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_711 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_735 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_754 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_788 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_800 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_859 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_915 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_941 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1057 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_478 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_540 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_690 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_700 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_761 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_827 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_887 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_319 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_380 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_440 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_560 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_618 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_668 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_752 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_786 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_803 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_859 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_915 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_947 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1057 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_148 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_247 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_580 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_772 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_778 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_887 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_943 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_957 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_963 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_975 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_987 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_170 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_400 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_555 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_808 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_842 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_848 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_915 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_965 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1057 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_296 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_342 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_548 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_640 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_696 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_791 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_812 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_871 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_883 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_943 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_975 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_554 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_600 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_621 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_650 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_731 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_831 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_844 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_915 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_971 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_985 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_991 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1003 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1015 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1057 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_124 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_198 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_353 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_400 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_467 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_612 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_660 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_772 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_827 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_857 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_886 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_943 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_975 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_993 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_315 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_325 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_575 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_582 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_780 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_786 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_833 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_846 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_854 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_899 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_911 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_971 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_997 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1003 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1015 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1052 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1058 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_148 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_355 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_466 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_774 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_796 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_830 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_864 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_943 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_975 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_999 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1013 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1025 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_315 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_462 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_719 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_836 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_840 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_862 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_888 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_971 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1003 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1015 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1047 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_124 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_189 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_310 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_478 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_543 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_646 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_659 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_703 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_716 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_886 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_943 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_975 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_999 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1031 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1055 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_90 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_504 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_526 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_568 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_650 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_715 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_743 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_800 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_806 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_834 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_840 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_846 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_852 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_862 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_915 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_971 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1003 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1027 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1041 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1057 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_128 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_300 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_409 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_476 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_692 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_711 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_740 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_760 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_790 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_882 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_943 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_975 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_999 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1031 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1055 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_106 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_260 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_388 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_443 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_668 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_712 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_718 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_786 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_822 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_844 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_874 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_878 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_971 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1003 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1027 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1047 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1053 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_267 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_301 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_386 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_488 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_572 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_628 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_747 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_920 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_926 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_932 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_938 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_975 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_999 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1031 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1055 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_490 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_728 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_802 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_832 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_855 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_874 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_971 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1003 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1027 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1047 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_134 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_348 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_366 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_595 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_770 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_846 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_874 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_943 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_975 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_999 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1031 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_448 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_620 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_730 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_817 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_898 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_904 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_910 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_971 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1003 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1027 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1047 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1053 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_528 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_662 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_707 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_836 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_854 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_886 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_943 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_975 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_999 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1031 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1055 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_270 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_384 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_456 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_509 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_576 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_640 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_712 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_840 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_878 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_888 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_915 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_971 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1003 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1027 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_1041 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1052 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1058 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_92 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_191 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_354 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_522 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_528 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_703 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_774 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_943 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_975 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_999 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1031 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1043 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1052 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_103 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_322 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_440 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_528 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_556 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_563 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_658 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_767 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_788 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_836 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_849 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_855 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_899 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_911 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_971 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1003 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1027 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_1044 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1052 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1057 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_523 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_634 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_679 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_683 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_733 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_838 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_876 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_882 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_943 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_975 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_999 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1019 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1025 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1031 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1044 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_100 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_172 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_269 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_340 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_431 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_663 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_676 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_788 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_802 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_824 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_874 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_886 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_892 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_898 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_904 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_910 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_971 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1003 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1015 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1044 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1053 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_71 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_252 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_428 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_480 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_509 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_747 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_760 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_807 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_861 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_887 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_943 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_975 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_999 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1025 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_1031 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1044 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1048 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1052 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1058 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_120 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_283 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_340 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_575 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_684 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_724 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_796 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_886 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_892 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_898 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_904 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_910 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_971 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1003 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1027 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_1041 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1052 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1058 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_70 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_187 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_406 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_486 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_518 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_871 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_886 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_943 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_975 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_999 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1025 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_443 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_514 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_568 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_659 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_665 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_800 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_848 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_854 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_892 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_898 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_904 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_910 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_971 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1003 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1027 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1047 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1053 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_131 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_264 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_274 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_411 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_800 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_827 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_846 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_927 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_939 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_975 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_999 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1031 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1055 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_70 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_259 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_456 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_578 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_856 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_900 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_912 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_971 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1003 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1027 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1047 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1053 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_66 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_127 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_368 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_532 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_874 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_883 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_943 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_975 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_999 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1031 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1055 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_275 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_358 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_388 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_768 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_836 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_911 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_971 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1003 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1027 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1041 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_67 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_148 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_245 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_478 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_565 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_756 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_795 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_831 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_837 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_873 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_920 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_926 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_932 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_938 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_975 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_999 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1031 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1055 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_323 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_435 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_665 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_746 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_779 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_900 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_912 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_971 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1003 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1027 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1047 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1053 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_355 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_444 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_518 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_694 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_704 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_750 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_762 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_790 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_828 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_859 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_868 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_943 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_975 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_999 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1031 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1055 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_378 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_600 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_674 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_722 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_728 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_788 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_810 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_836 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_858 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_899 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_911 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_971 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1003 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1027 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1047 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1053 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_86 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_245 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_398 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_467 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_566 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_588 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_734 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_767 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_789 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_864 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_943 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_975 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_999 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1031 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_227 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_672 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_834 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_900 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_912 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_971 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1003 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1027 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1047 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_72 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_259 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_690 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_747 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_801 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_859 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_872 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_943 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_975 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_999 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1031 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1055 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_314 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_327 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_686 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_730 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_779 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_824 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_852 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_882 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_889 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_971 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1003 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1027 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1047 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1053 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_131 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_191 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_357 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_556 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_780 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_864 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_871 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_878 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_887 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_943 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_975 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_999 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1031 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1055 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_94 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_448 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_516 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_596 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_746 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_831 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_856 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_899 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_911 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_971 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1003 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1027 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1041 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1057 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_424 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_516 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_546 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_582 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_628 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_652 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_770 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_796 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_816 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_846 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_870 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_943 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_975 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_999 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1031 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1052 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_215 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_336 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_392 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_512 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_548 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_556 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_778 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_840 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_900 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_912 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_971 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1003 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1027 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_1041 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_1052 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1058 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_758 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_806 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_872 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_943 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_975 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_999 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1031 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1055 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_466 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_551 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_656 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_752 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_806 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_827 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_840 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_846 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_890 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_971 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1003 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1027 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1047 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_1053 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_534 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_703 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_768 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_781 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_854 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_902 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_975 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_999 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1031 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_269 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_385 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_548 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_560 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_568 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_683 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_799 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_806 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_866 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_896 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_971 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1003 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1027 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1047 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_1053 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_130 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_316 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_467 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_628 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_656 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_691 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_703 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_801 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_864 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_872 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_920 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_926 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_932 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_938 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_975 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_999 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1031 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1055 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_71 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_158 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_344 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_439 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_656 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_781 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_899 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_911 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_971 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1003 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1027 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1047 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_1053 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_61 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_87 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_182 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_348 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_510 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_726 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_866 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_870 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_880 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_943 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_975 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_999 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1031 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1055 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_728 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_732 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_859 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_971 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1003 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1027 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1041 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1057 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_200 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_592 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_702 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_830 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_882 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_943 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_975 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_999 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1031 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1043 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1052 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1058 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_134 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_344 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_439 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_516 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_526 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_786 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_840 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_898 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_904 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_910 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_971 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1003 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1027 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1047 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_75 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_357 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_509 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_686 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_799 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_816 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_864 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_872 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_928 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_934 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_940 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_975 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_999 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1031 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1055 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_497 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_674 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_743 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_779 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_866 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_878 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_898 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_911 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_971 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1003 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1027 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1047 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_1053 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_399 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_538 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_572 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_628 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_644 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_700 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_804 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_846 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_854 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_912 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_927 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_939 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_975 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_999 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1031 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_78 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_607 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_640 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_677 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_731 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_792 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_842 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_866 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_882 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_892 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_898 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_904 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_910 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_971 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1003 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1027 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1047 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1053 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_267 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_303 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_372 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_411 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_544 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_581 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_628 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_691 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_845 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_851 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_861 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_880 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_943 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_975 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_999 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1031 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1055 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_504 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_728 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_831 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_846 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_889 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_915 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_971 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1003 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1027 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1047 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_300 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_470 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_648 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_693 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_768 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_793 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_838 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_883 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_920 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_926 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_932 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_938 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_975 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_999 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1031 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1055 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_466 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_515 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_622 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_660 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_696 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_720 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_730 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_746 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_817 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_854 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_874 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_898 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_911 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_971 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1003 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1027 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1041 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1057 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_130 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_350 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_481 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_510 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_603 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_646 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_691 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_796 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_864 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_872 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_894 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_911 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_920 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_926 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_932 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_938 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_975 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_999 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1031 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_1043 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_1052 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1058 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_40 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_327 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_619 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_684 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_843 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_866 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_910 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_971 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1003 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1027 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1047 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_75 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_118 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_528 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_579 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_697 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_739 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_943 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_975 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_999 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1031 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1055 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_56 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_227 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_426 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_452 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_516 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_624 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_789 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_825 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_847 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_874 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_971 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1003 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1027 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1047 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_1053 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_191 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_370 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_511 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_684 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_714 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_771 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_883 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_887 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_916 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_928 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_934 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_940 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_975 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_999 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1031 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_58 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_103 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_444 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_631 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_732 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_818 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_843 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_876 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_898 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_915 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_971 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1003 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1027 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1047 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1053 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_187 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_191 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_254 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_357 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_846 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_878 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_943 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_975 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_999 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1031 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1055 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_47 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_64 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_179 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_344 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_439 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_624 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_656 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_851 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_890 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_915 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_971 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1003 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1027 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1047 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_40 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_61 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_295 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_316 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_634 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_827 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_859 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_943 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_975 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_999 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1031 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1055 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_215 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_274 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_325 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_552 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_663 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_676 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_775 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_858 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_911 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_971 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1003 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1027 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1041 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_30 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_75 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_106 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_539 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_566 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_684 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_920 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_926 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_932 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_938 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_975 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_999 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1031 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1055 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_383 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_516 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_568 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_690 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_724 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_806 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_892 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_912 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_971 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1003 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1027 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1047 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_1053 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_127 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_245 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_424 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_638 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_790 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_812 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_818 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_828 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_852 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_876 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_920 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_926 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_932 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_938 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_975 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_999 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1031 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1055 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_259 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_508 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_578 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_656 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_677 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_714 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_799 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_811 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_832 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_858 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_886 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_892 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_898 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_904 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_910 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_971 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1003 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1027 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1047 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_424 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_537 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_652 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_678 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_887 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_943 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_975 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_999 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1031 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_226 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_512 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_552 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_600 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_668 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_674 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_786 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_798 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_834 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_848 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_855 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_888 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_971 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_1003 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_1027 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_1047 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_1053 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_40 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_124 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_372 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_536 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_588 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_602 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_621 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_652 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_695 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_702 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_864 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_884 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_943 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_975 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_999 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1031 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1055 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_159 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_344 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_396 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_450 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_519 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_650 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_680 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_786 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_806 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_854 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_878 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_884 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_890 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_896 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_971 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_1003 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_1027 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_244 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_299 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_312 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_579 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_621 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_678 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_816 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_830 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_855 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_867 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_886 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_943 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_975 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_999 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1013 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1019 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1031 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1055 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_228 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_382 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_551 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_612 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_667 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_717 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_788 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_834 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_840 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_844 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_854 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_876 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_882 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_888 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_892 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_896 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_971 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_1003 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1015 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_135 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_398 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_540 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_604 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_772 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_815 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_887 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_943 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_975 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_999 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_99 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_315 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_638 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_672 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_817 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_899 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_911 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_971 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_991 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_997 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1057 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_635 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_648 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_747 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_754 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_865 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_943 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_975 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_987 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_98 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_343 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_526 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_672 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_798 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_848 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_874 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_886 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_892 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_898 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_904 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_910 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_971 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1057 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_124 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_413 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_491 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_571 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_646 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_700 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_733 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_772 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_802 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_814 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_818 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_824 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_856 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_862 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_883 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_920 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_926 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_932 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_938 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_963 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_969 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_275 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_384 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_509 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_555 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_599 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_656 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_674 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_697 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_707 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_752 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_779 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_803 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_855 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_915 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_971 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1057 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_135 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_142 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_677 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_705 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_751 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_796 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_836 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_943 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_963 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_969 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_158 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_519 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_602 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_742 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_762 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_831 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_844 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_899 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_911 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_971 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1057 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_131 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_366 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_602 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_760 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_789 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_806 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_874 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_887 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_943 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_969 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_975 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_987 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_102 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_395 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_539 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_723 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_788 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_824 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_830 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_836 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_846 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_915 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_971 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_1057 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_187 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_245 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_536 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_635 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_648 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_772 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_808 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_814 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_838 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_862 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_868 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_874 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_886 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_943 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_963 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_969 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_684 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_796 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_818 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_879 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_900 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_912 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_965 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_1057 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_378 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_526 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_595 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_679 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_771 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_778 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_871 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_884 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_943 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_957 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_963 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_975 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_987 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_114 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_578 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_707 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_731 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_878 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_884 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_890 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_896 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_947 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_1057 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_118 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_355 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_524 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_760 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_764 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_801 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_805 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_852 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_858 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_866 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_874 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_887 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_920 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_926 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_932 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_938 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_146 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_172 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_385 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_444 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_560 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_599 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_674 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_783 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_859 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_915 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_959 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_342 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_404 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_544 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_627 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_683 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_748 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_828 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_887 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_943 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_400 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_499 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_568 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_654 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_783 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_836 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_842 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_848 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_854 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_915 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_935 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_941 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_1057 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_484 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_588 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_640 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_650 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_700 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_828 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_887 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_931 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_147 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_515 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_526 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_728 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_742 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_859 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_915 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_941 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_1057 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_179 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_288 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_316 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_420 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_484 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_566 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_658 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_700 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_745 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_758 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_806 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_836 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_848 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_854 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_872 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_878 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_884 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_919 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_623 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_803 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_859 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_915 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_941 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_344 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_366 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_467 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_636 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_738 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_758 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_808 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_814 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_887 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_931 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_336 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_548 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_632 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_665 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_728 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_834 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_840 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_846 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_915 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_935 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_947 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_959 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_1057 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_182 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_357 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_423 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_463 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_546 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_659 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_770 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_814 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_820 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_848 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_854 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_872 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_878 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_884 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_931 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_154 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_400 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_454 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_574 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_616 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_624 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_716 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_778 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_799 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_859 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_915 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_941 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_947 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_959 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1057 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_259 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_311 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_355 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_512 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_547 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_582 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_622 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_634 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_677 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_767 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_800 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_806 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_814 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_887 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_176 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_560 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_672 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_799 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_833 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_843 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_915 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_941 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_947 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_959 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_1057 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_74 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_322 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_368 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_704 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_749 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_756 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_794 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_855 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_861 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_943 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_163 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_288 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_560 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_623 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_665 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_674 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_731 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_774 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_803 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_847 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_855 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_915 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_947 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_230 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_626 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_677 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_702 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_756 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_767 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_800 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_806 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_848 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_854 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_872 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_878 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_884 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_943 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_957 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_969 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_215 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_344 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_395 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_537 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_660 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_748 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_773 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_846 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_915 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_941 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_947 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_959 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_1057 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_30 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_34 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_140 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_466 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_550 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_606 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_705 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_756 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_830 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_871 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_883 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_943 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_957 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_969 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_316 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_498 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_515 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_575 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_640 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_742 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_766 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_828 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_843 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_854 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_915 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_959 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_548 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_660 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_684 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_848 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_854 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_872 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_878 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_884 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_911 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_917 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_957 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_969 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1057 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_282 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_542 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_560 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_572 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_582 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_664 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_731 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_786 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_915 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_947 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_235 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_574 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_696 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_791 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_851 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_857 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_870 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_876 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_882 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_943 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1057 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_78 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_329 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_539 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_640 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_658 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_788 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_799 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_806 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_843 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_855 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_915 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_935 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_947 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_959 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_19 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_72 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_357 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_366 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_428 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_480 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_583 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_591 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_637 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_799 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_806 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_887 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_931 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1057 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_459 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_556 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_600 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_656 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_665 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_731 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_767 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_859 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_915 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_1057 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_17 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_202 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_427 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_599 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_683 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_703 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_756 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_887 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_907 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_913 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_466 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_495 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_636 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_786 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_859 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_903 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_316 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_352 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_372 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_546 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_658 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_696 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_748 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_836 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_848 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_854 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_872 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_878 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_884 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_901 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_913 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_94 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_179 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_264 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_553 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_675 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_733 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_802 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_859 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_885 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_891 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_13 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_67 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_242 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_308 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_459 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_548 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_762 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_814 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_887 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_16 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_25 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_48 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_215 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_343 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_437 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_466 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_508 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_599 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_631 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_638 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_658 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_674 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_715 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_859 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_879 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_885 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_87 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_355 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_364 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_470 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_511 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_736 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_760 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_828 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_875 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_46 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_387 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_438 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_560 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_606 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_723 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_773 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_800 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_835 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_885 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_891 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_230 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_480 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_602 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_610 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_668 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_693 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_700 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_881 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_24 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_459 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_551 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_655 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_664 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_728 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_803 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_859 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_879 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_885 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_13 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_30 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_476 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_628 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_677 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_724 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_758 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_773 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_806 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_831 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_875 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1057 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_49 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_70 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_155 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_219 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_550 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_640 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_663 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_674 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_724 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_836 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_842 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_848 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_854 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_873 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_879 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_891 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_1057 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_256 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_547 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_658 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_703 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_747 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_763 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_814 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_881 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1057 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_48 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_126 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_284 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_507 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_511 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_560 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_728 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_859 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_885 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_891 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_1057 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_84 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_260 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_367 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_467 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_527 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_628 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_655 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_708 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_743 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_827 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_875 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_103 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_134 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_487 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_507 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_560 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_582 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_624 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_717 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_767 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_859 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_873 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_879 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_891 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_319 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_330 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_431 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_572 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_644 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_654 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_771 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_807 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1057 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_114 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_228 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_259 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_292 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_327 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_508 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_572 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_666 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_716 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_740 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_859 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_322 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_413 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_484 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_522 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_679 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_700 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_771 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_831 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_851 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_857 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_215 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_504 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_539 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_575 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_634 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_661 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_723 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_803 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_847 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_135 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_191 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_288 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_470 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_478 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_658 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_700 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_708 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_758 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_831 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_857 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_100 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_179 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_435 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_521 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_616 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_623 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_667 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_680 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_720 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_730 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_803 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_829 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_835 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_847 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_592 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_633 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_697 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_825 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_846 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_858 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_870 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_146 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_315 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_387 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_494 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_509 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_735 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_786 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_823 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_829 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_142 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_428 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_494 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_603 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_628 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_652 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_819 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_394 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_452 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_456 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_494 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_537 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_627 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_660 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_803 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_817 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_829 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_42 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_186 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_372 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_398 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_588 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_703 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_459 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_470 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_576 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_593 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_631 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_651 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_668 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_716 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_787 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_799 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_817 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_829 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_1057 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_183 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_366 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_490 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_638 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_660 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_666 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_807 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_235 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_370 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_450 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_560 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_607 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_624 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_791 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_1057 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_140 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_330 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_343 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_480 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_595 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_758 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_795 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_807 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_269 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_494 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_518 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_544 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_575 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_667 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_719 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_779 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_1057 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_479 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_600 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_171 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_404 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_515 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_604 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_740 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_767 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_779 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_1057 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_353 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_378 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_466 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_516 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_547 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_758 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_396 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_537 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_554 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_560 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_1057 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_332 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_410 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_483 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_495 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_526 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_543 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_580 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_604 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_633 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_703 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_715 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_739 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_406 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_544 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_603 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_330 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_439 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_578 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_470 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_535 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_495 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_550 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_723 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_434 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_470 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_528 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_540 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_580 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_689 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_749 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_771 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1033 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_580 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_745 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_818 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_848 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_860 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_986 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1014 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1034 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_1046 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1052 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1057 ();
 assign mem_addr[24] = net98;
 assign mem_addr[25] = net99;
 assign mem_addr[26] = net100;
 assign mem_addr[27] = net101;
 assign mem_addr[28] = net102;
 assign mem_addr[29] = net103;
 assign mem_addr[30] = net104;
 assign mem_addr[31] = net105;
endmodule

